** Cell name: sram_64x4
.subckt sram_64x4 vdd gnd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] in_b[0] in_b[1] in_b[2] in_b[3] in_b[4] in_b[5] in_b[6] in_b[7] in_b[8] in_b[9] in_b[10] in_b[11] in_b[12] in_b[13] in_b[14] in_b[15] in_b[16] in_b[17] in_b[18] in_b[19] in_b[20] in_b[21] in_b[22] in_b[23] in_b[24] in_b[25] in_b[26] in_b[27] in_b[28] in_b[29] in_b[30] in_b[31] in_b[32] in_b[33] in_b[34] in_b[35] in_b[36] in_b[37] in_b[38] in_b[39] in_b[40] in_b[41] in_b[42] in_b[43] in_b[44] in_b[45] in_b[46] in_b[47] in_b[48] in_b[49] in_b[50] in_b[51] in_b[52] in_b[53] in_b[54] in_b[55] in_b[56] in_b[57] in_b[58] in_b[59] in_b[60] in_b[61] in_b[62] in_b[63] bl[0] bl[1] bl[2] bl[3] bl_b[0] bl_b[1] bl_b[2] bl_b[3] bitcell_out_0[0] bitcell_out_0[1] bitcell_out_0[2] bitcell_out_0[3] bitcell_out_1[0] bitcell_out_1[1] bitcell_out_1[2] bitcell_out_1[3] bitcell_out_2[0] bitcell_out_2[1] bitcell_out_2[2] bitcell_out_2[3] bitcell_out_3[0] bitcell_out_3[1] bitcell_out_3[2] bitcell_out_3[3] bitcell_out_4[0] bitcell_out_4[1] bitcell_out_4[2] bitcell_out_4[3] bitcell_out_5[0] bitcell_out_5[1] bitcell_out_5[2] bitcell_out_5[3] bitcell_out_6[0] bitcell_out_6[1] bitcell_out_6[2] bitcell_out_6[3] bitcell_out_7[0] bitcell_out_7[1] bitcell_out_7[2] bitcell_out_7[3] bitcell_out_8[0] bitcell_out_8[1] bitcell_out_8[2] bitcell_out_8[3] bitcell_out_9[0] bitcell_out_9[1] bitcell_out_9[2] bitcell_out_9[3] bitcell_out_10[0] bitcell_out_10[1] bitcell_out_10[2] bitcell_out_10[3] bitcell_out_11[0] bitcell_out_11[1] bitcell_out_11[2] bitcell_out_11[3] bitcell_out_12[0] bitcell_out_12[1] bitcell_out_12[2] bitcell_out_12[3] bitcell_out_13[0] bitcell_out_13[1] bitcell_out_13[2] bitcell_out_13[3] bitcell_out_14[0] bitcell_out_14[1] bitcell_out_14[2] bitcell_out_14[3] bitcell_out_15[0] bitcell_out_15[1] bitcell_out_15[2] bitcell_out_15[3] bitcell_out_16[0] bitcell_out_16[1] bitcell_out_16[2] bitcell_out_16[3] bitcell_out_17[0] bitcell_out_17[1] bitcell_out_17[2] bitcell_out_17[3] bitcell_out_18[0] bitcell_out_18[1] bitcell_out_18[2] bitcell_out_18[3] bitcell_out_19[0] bitcell_out_19[1] bitcell_out_19[2] bitcell_out_19[3] bitcell_out_20[0] bitcell_out_20[1] bitcell_out_20[2] bitcell_out_20[3] bitcell_out_21[0] bitcell_out_21[1] bitcell_out_21[2] bitcell_out_21[3] bitcell_out_22[0] bitcell_out_22[1] bitcell_out_22[2] bitcell_out_22[3] bitcell_out_23[0] bitcell_out_23[1] bitcell_out_23[2] bitcell_out_23[3] bitcell_out_24[0] bitcell_out_24[1] bitcell_out_24[2] bitcell_out_24[3] bitcell_out_25[0] bitcell_out_25[1] bitcell_out_25[2] bitcell_out_25[3] bitcell_out_26[0] bitcell_out_26[1] bitcell_out_26[2] bitcell_out_26[3] bitcell_out_27[0] bitcell_out_27[1] bitcell_out_27[2] bitcell_out_27[3] bitcell_out_28[0] bitcell_out_28[1] bitcell_out_28[2] bitcell_out_28[3] bitcell_out_29[0] bitcell_out_29[1] bitcell_out_29[2] bitcell_out_29[3] bitcell_out_30[0] bitcell_out_30[1] bitcell_out_30[2] bitcell_out_30[3] bitcell_out_31[0] bitcell_out_31[1] bitcell_out_31[2] bitcell_out_31[3] bitcell_out_32[0] bitcell_out_32[1] bitcell_out_32[2] bitcell_out_32[3] bitcell_out_33[0] bitcell_out_33[1] bitcell_out_33[2] bitcell_out_33[3] bitcell_out_34[0] bitcell_out_34[1] bitcell_out_34[2] bitcell_out_34[3] bitcell_out_35[0] bitcell_out_35[1] bitcell_out_35[2] bitcell_out_35[3] bitcell_out_36[0] bitcell_out_36[1] bitcell_out_36[2] bitcell_out_36[3] bitcell_out_37[0] bitcell_out_37[1] bitcell_out_37[2] bitcell_out_37[3] bitcell_out_38[0] bitcell_out_38[1] bitcell_out_38[2] bitcell_out_38[3] bitcell_out_39[0] bitcell_out_39[1] bitcell_out_39[2] bitcell_out_39[3] bitcell_out_40[0] bitcell_out_40[1] bitcell_out_40[2] bitcell_out_40[3] bitcell_out_41[0] bitcell_out_41[1] bitcell_out_41[2] bitcell_out_41[3] bitcell_out_42[0] bitcell_out_42[1] bitcell_out_42[2] bitcell_out_42[3] bitcell_out_43[0] bitcell_out_43[1] bitcell_out_43[2] bitcell_out_43[3] bitcell_out_44[0] bitcell_out_44[1] bitcell_out_44[2] bitcell_out_44[3] bitcell_out_45[0] bitcell_out_45[1] bitcell_out_45[2] bitcell_out_45[3] bitcell_out_46[0] bitcell_out_46[1] bitcell_out_46[2] bitcell_out_46[3] bitcell_out_47[0] bitcell_out_47[1] bitcell_out_47[2] bitcell_out_47[3] bitcell_out_48[0] bitcell_out_48[1] bitcell_out_48[2] bitcell_out_48[3] bitcell_out_49[0] bitcell_out_49[1] bitcell_out_49[2] bitcell_out_49[3] bitcell_out_50[0] bitcell_out_50[1] bitcell_out_50[2] bitcell_out_50[3] bitcell_out_51[0] bitcell_out_51[1] bitcell_out_51[2] bitcell_out_51[3] bitcell_out_52[0] bitcell_out_52[1] bitcell_out_52[2] bitcell_out_52[3] bitcell_out_53[0] bitcell_out_53[1] bitcell_out_53[2] bitcell_out_53[3] bitcell_out_54[0] bitcell_out_54[1] bitcell_out_54[2] bitcell_out_54[3] bitcell_out_55[0] bitcell_out_55[1] bitcell_out_55[2] bitcell_out_55[3] bitcell_out_56[0] bitcell_out_56[1] bitcell_out_56[2] bitcell_out_56[3] bitcell_out_57[0] bitcell_out_57[1] bitcell_out_57[2] bitcell_out_57[3] bitcell_out_58[0] bitcell_out_58[1] bitcell_out_58[2] bitcell_out_58[3] bitcell_out_59[0] bitcell_out_59[1] bitcell_out_59[2] bitcell_out_59[3] bitcell_out_60[0] bitcell_out_60[1] bitcell_out_60[2] bitcell_out_60[3] bitcell_out_61[0] bitcell_out_61[1] bitcell_out_61[2] bitcell_out_61[3] bitcell_out_62[0] bitcell_out_62[1] bitcell_out_62[2] bitcell_out_62[3] bitcell_out_63[0] bitcell_out_63[1] bitcell_out_63[2] bitcell_out_63[3] 
xi_bitcell_0_0 vdd gnd wl[0] in_b[0] bl[0] bl_b[0] bitcell_out_0[0] dcim_bitcell
xi_bitcell_0_1 vdd gnd wl[0] in_b[0] bl[1] bl_b[1] bitcell_out_0[1] dcim_bitcell
xi_bitcell_0_2 vdd gnd wl[0] in_b[0] bl[2] bl_b[2] bitcell_out_0[2] dcim_bitcell
xi_bitcell_0_3 vdd gnd wl[0] in_b[0] bl[3] bl_b[3] bitcell_out_0[3] dcim_bitcell
xi_bitcell_1_0 vdd gnd wl[1] in_b[1] bl[0] bl_b[0] bitcell_out_1[0] dcim_bitcell
xi_bitcell_1_1 vdd gnd wl[1] in_b[1] bl[1] bl_b[1] bitcell_out_1[1] dcim_bitcell
xi_bitcell_1_2 vdd gnd wl[1] in_b[1] bl[2] bl_b[2] bitcell_out_1[2] dcim_bitcell
xi_bitcell_1_3 vdd gnd wl[1] in_b[1] bl[3] bl_b[3] bitcell_out_1[3] dcim_bitcell
xi_bitcell_2_0 vdd gnd wl[2] in_b[2] bl[0] bl_b[0] bitcell_out_2[0] dcim_bitcell
xi_bitcell_2_1 vdd gnd wl[2] in_b[2] bl[1] bl_b[1] bitcell_out_2[1] dcim_bitcell
xi_bitcell_2_2 vdd gnd wl[2] in_b[2] bl[2] bl_b[2] bitcell_out_2[2] dcim_bitcell
xi_bitcell_2_3 vdd gnd wl[2] in_b[2] bl[3] bl_b[3] bitcell_out_2[3] dcim_bitcell
xi_bitcell_3_0 vdd gnd wl[3] in_b[3] bl[0] bl_b[0] bitcell_out_3[0] dcim_bitcell
xi_bitcell_3_1 vdd gnd wl[3] in_b[3] bl[1] bl_b[1] bitcell_out_3[1] dcim_bitcell
xi_bitcell_3_2 vdd gnd wl[3] in_b[3] bl[2] bl_b[2] bitcell_out_3[2] dcim_bitcell
xi_bitcell_3_3 vdd gnd wl[3] in_b[3] bl[3] bl_b[3] bitcell_out_3[3] dcim_bitcell
xi_bitcell_4_0 vdd gnd wl[4] in_b[4] bl[0] bl_b[0] bitcell_out_4[0] dcim_bitcell
xi_bitcell_4_1 vdd gnd wl[4] in_b[4] bl[1] bl_b[1] bitcell_out_4[1] dcim_bitcell
xi_bitcell_4_2 vdd gnd wl[4] in_b[4] bl[2] bl_b[2] bitcell_out_4[2] dcim_bitcell
xi_bitcell_4_3 vdd gnd wl[4] in_b[4] bl[3] bl_b[3] bitcell_out_4[3] dcim_bitcell
xi_bitcell_5_0 vdd gnd wl[5] in_b[5] bl[0] bl_b[0] bitcell_out_5[0] dcim_bitcell
xi_bitcell_5_1 vdd gnd wl[5] in_b[5] bl[1] bl_b[1] bitcell_out_5[1] dcim_bitcell
xi_bitcell_5_2 vdd gnd wl[5] in_b[5] bl[2] bl_b[2] bitcell_out_5[2] dcim_bitcell
xi_bitcell_5_3 vdd gnd wl[5] in_b[5] bl[3] bl_b[3] bitcell_out_5[3] dcim_bitcell
xi_bitcell_6_0 vdd gnd wl[6] in_b[6] bl[0] bl_b[0] bitcell_out_6[0] dcim_bitcell
xi_bitcell_6_1 vdd gnd wl[6] in_b[6] bl[1] bl_b[1] bitcell_out_6[1] dcim_bitcell
xi_bitcell_6_2 vdd gnd wl[6] in_b[6] bl[2] bl_b[2] bitcell_out_6[2] dcim_bitcell
xi_bitcell_6_3 vdd gnd wl[6] in_b[6] bl[3] bl_b[3] bitcell_out_6[3] dcim_bitcell
xi_bitcell_7_0 vdd gnd wl[7] in_b[7] bl[0] bl_b[0] bitcell_out_7[0] dcim_bitcell
xi_bitcell_7_1 vdd gnd wl[7] in_b[7] bl[1] bl_b[1] bitcell_out_7[1] dcim_bitcell
xi_bitcell_7_2 vdd gnd wl[7] in_b[7] bl[2] bl_b[2] bitcell_out_7[2] dcim_bitcell
xi_bitcell_7_3 vdd gnd wl[7] in_b[7] bl[3] bl_b[3] bitcell_out_7[3] dcim_bitcell
xi_bitcell_8_0 vdd gnd wl[8] in_b[8] bl[0] bl_b[0] bitcell_out_8[0] dcim_bitcell
xi_bitcell_8_1 vdd gnd wl[8] in_b[8] bl[1] bl_b[1] bitcell_out_8[1] dcim_bitcell
xi_bitcell_8_2 vdd gnd wl[8] in_b[8] bl[2] bl_b[2] bitcell_out_8[2] dcim_bitcell
xi_bitcell_8_3 vdd gnd wl[8] in_b[8] bl[3] bl_b[3] bitcell_out_8[3] dcim_bitcell
xi_bitcell_9_0 vdd gnd wl[9] in_b[9] bl[0] bl_b[0] bitcell_out_9[0] dcim_bitcell
xi_bitcell_9_1 vdd gnd wl[9] in_b[9] bl[1] bl_b[1] bitcell_out_9[1] dcim_bitcell
xi_bitcell_9_2 vdd gnd wl[9] in_b[9] bl[2] bl_b[2] bitcell_out_9[2] dcim_bitcell
xi_bitcell_9_3 vdd gnd wl[9] in_b[9] bl[3] bl_b[3] bitcell_out_9[3] dcim_bitcell
xi_bitcell_10_0 vdd gnd wl[10] in_b[10] bl[0] bl_b[0] bitcell_out_10[0] dcim_bitcell
xi_bitcell_10_1 vdd gnd wl[10] in_b[10] bl[1] bl_b[1] bitcell_out_10[1] dcim_bitcell
xi_bitcell_10_2 vdd gnd wl[10] in_b[10] bl[2] bl_b[2] bitcell_out_10[2] dcim_bitcell
xi_bitcell_10_3 vdd gnd wl[10] in_b[10] bl[3] bl_b[3] bitcell_out_10[3] dcim_bitcell
xi_bitcell_11_0 vdd gnd wl[11] in_b[11] bl[0] bl_b[0] bitcell_out_11[0] dcim_bitcell
xi_bitcell_11_1 vdd gnd wl[11] in_b[11] bl[1] bl_b[1] bitcell_out_11[1] dcim_bitcell
xi_bitcell_11_2 vdd gnd wl[11] in_b[11] bl[2] bl_b[2] bitcell_out_11[2] dcim_bitcell
xi_bitcell_11_3 vdd gnd wl[11] in_b[11] bl[3] bl_b[3] bitcell_out_11[3] dcim_bitcell
xi_bitcell_12_0 vdd gnd wl[12] in_b[12] bl[0] bl_b[0] bitcell_out_12[0] dcim_bitcell
xi_bitcell_12_1 vdd gnd wl[12] in_b[12] bl[1] bl_b[1] bitcell_out_12[1] dcim_bitcell
xi_bitcell_12_2 vdd gnd wl[12] in_b[12] bl[2] bl_b[2] bitcell_out_12[2] dcim_bitcell
xi_bitcell_12_3 vdd gnd wl[12] in_b[12] bl[3] bl_b[3] bitcell_out_12[3] dcim_bitcell
xi_bitcell_13_0 vdd gnd wl[13] in_b[13] bl[0] bl_b[0] bitcell_out_13[0] dcim_bitcell
xi_bitcell_13_1 vdd gnd wl[13] in_b[13] bl[1] bl_b[1] bitcell_out_13[1] dcim_bitcell
xi_bitcell_13_2 vdd gnd wl[13] in_b[13] bl[2] bl_b[2] bitcell_out_13[2] dcim_bitcell
xi_bitcell_13_3 vdd gnd wl[13] in_b[13] bl[3] bl_b[3] bitcell_out_13[3] dcim_bitcell
xi_bitcell_14_0 vdd gnd wl[14] in_b[14] bl[0] bl_b[0] bitcell_out_14[0] dcim_bitcell
xi_bitcell_14_1 vdd gnd wl[14] in_b[14] bl[1] bl_b[1] bitcell_out_14[1] dcim_bitcell
xi_bitcell_14_2 vdd gnd wl[14] in_b[14] bl[2] bl_b[2] bitcell_out_14[2] dcim_bitcell
xi_bitcell_14_3 vdd gnd wl[14] in_b[14] bl[3] bl_b[3] bitcell_out_14[3] dcim_bitcell
xi_bitcell_15_0 vdd gnd wl[15] in_b[15] bl[0] bl_b[0] bitcell_out_15[0] dcim_bitcell
xi_bitcell_15_1 vdd gnd wl[15] in_b[15] bl[1] bl_b[1] bitcell_out_15[1] dcim_bitcell
xi_bitcell_15_2 vdd gnd wl[15] in_b[15] bl[2] bl_b[2] bitcell_out_15[2] dcim_bitcell
xi_bitcell_15_3 vdd gnd wl[15] in_b[15] bl[3] bl_b[3] bitcell_out_15[3] dcim_bitcell
xi_bitcell_16_0 vdd gnd wl[16] in_b[16] bl[0] bl_b[0] bitcell_out_16[0] dcim_bitcell
xi_bitcell_16_1 vdd gnd wl[16] in_b[16] bl[1] bl_b[1] bitcell_out_16[1] dcim_bitcell
xi_bitcell_16_2 vdd gnd wl[16] in_b[16] bl[2] bl_b[2] bitcell_out_16[2] dcim_bitcell
xi_bitcell_16_3 vdd gnd wl[16] in_b[16] bl[3] bl_b[3] bitcell_out_16[3] dcim_bitcell
xi_bitcell_17_0 vdd gnd wl[17] in_b[17] bl[0] bl_b[0] bitcell_out_17[0] dcim_bitcell
xi_bitcell_17_1 vdd gnd wl[17] in_b[17] bl[1] bl_b[1] bitcell_out_17[1] dcim_bitcell
xi_bitcell_17_2 vdd gnd wl[17] in_b[17] bl[2] bl_b[2] bitcell_out_17[2] dcim_bitcell
xi_bitcell_17_3 vdd gnd wl[17] in_b[17] bl[3] bl_b[3] bitcell_out_17[3] dcim_bitcell
xi_bitcell_18_0 vdd gnd wl[18] in_b[18] bl[0] bl_b[0] bitcell_out_18[0] dcim_bitcell
xi_bitcell_18_1 vdd gnd wl[18] in_b[18] bl[1] bl_b[1] bitcell_out_18[1] dcim_bitcell
xi_bitcell_18_2 vdd gnd wl[18] in_b[18] bl[2] bl_b[2] bitcell_out_18[2] dcim_bitcell
xi_bitcell_18_3 vdd gnd wl[18] in_b[18] bl[3] bl_b[3] bitcell_out_18[3] dcim_bitcell
xi_bitcell_19_0 vdd gnd wl[19] in_b[19] bl[0] bl_b[0] bitcell_out_19[0] dcim_bitcell
xi_bitcell_19_1 vdd gnd wl[19] in_b[19] bl[1] bl_b[1] bitcell_out_19[1] dcim_bitcell
xi_bitcell_19_2 vdd gnd wl[19] in_b[19] bl[2] bl_b[2] bitcell_out_19[2] dcim_bitcell
xi_bitcell_19_3 vdd gnd wl[19] in_b[19] bl[3] bl_b[3] bitcell_out_19[3] dcim_bitcell
xi_bitcell_20_0 vdd gnd wl[20] in_b[20] bl[0] bl_b[0] bitcell_out_20[0] dcim_bitcell
xi_bitcell_20_1 vdd gnd wl[20] in_b[20] bl[1] bl_b[1] bitcell_out_20[1] dcim_bitcell
xi_bitcell_20_2 vdd gnd wl[20] in_b[20] bl[2] bl_b[2] bitcell_out_20[2] dcim_bitcell
xi_bitcell_20_3 vdd gnd wl[20] in_b[20] bl[3] bl_b[3] bitcell_out_20[3] dcim_bitcell
xi_bitcell_21_0 vdd gnd wl[21] in_b[21] bl[0] bl_b[0] bitcell_out_21[0] dcim_bitcell
xi_bitcell_21_1 vdd gnd wl[21] in_b[21] bl[1] bl_b[1] bitcell_out_21[1] dcim_bitcell
xi_bitcell_21_2 vdd gnd wl[21] in_b[21] bl[2] bl_b[2] bitcell_out_21[2] dcim_bitcell
xi_bitcell_21_3 vdd gnd wl[21] in_b[21] bl[3] bl_b[3] bitcell_out_21[3] dcim_bitcell
xi_bitcell_22_0 vdd gnd wl[22] in_b[22] bl[0] bl_b[0] bitcell_out_22[0] dcim_bitcell
xi_bitcell_22_1 vdd gnd wl[22] in_b[22] bl[1] bl_b[1] bitcell_out_22[1] dcim_bitcell
xi_bitcell_22_2 vdd gnd wl[22] in_b[22] bl[2] bl_b[2] bitcell_out_22[2] dcim_bitcell
xi_bitcell_22_3 vdd gnd wl[22] in_b[22] bl[3] bl_b[3] bitcell_out_22[3] dcim_bitcell
xi_bitcell_23_0 vdd gnd wl[23] in_b[23] bl[0] bl_b[0] bitcell_out_23[0] dcim_bitcell
xi_bitcell_23_1 vdd gnd wl[23] in_b[23] bl[1] bl_b[1] bitcell_out_23[1] dcim_bitcell
xi_bitcell_23_2 vdd gnd wl[23] in_b[23] bl[2] bl_b[2] bitcell_out_23[2] dcim_bitcell
xi_bitcell_23_3 vdd gnd wl[23] in_b[23] bl[3] bl_b[3] bitcell_out_23[3] dcim_bitcell
xi_bitcell_24_0 vdd gnd wl[24] in_b[24] bl[0] bl_b[0] bitcell_out_24[0] dcim_bitcell
xi_bitcell_24_1 vdd gnd wl[24] in_b[24] bl[1] bl_b[1] bitcell_out_24[1] dcim_bitcell
xi_bitcell_24_2 vdd gnd wl[24] in_b[24] bl[2] bl_b[2] bitcell_out_24[2] dcim_bitcell
xi_bitcell_24_3 vdd gnd wl[24] in_b[24] bl[3] bl_b[3] bitcell_out_24[3] dcim_bitcell
xi_bitcell_25_0 vdd gnd wl[25] in_b[25] bl[0] bl_b[0] bitcell_out_25[0] dcim_bitcell
xi_bitcell_25_1 vdd gnd wl[25] in_b[25] bl[1] bl_b[1] bitcell_out_25[1] dcim_bitcell
xi_bitcell_25_2 vdd gnd wl[25] in_b[25] bl[2] bl_b[2] bitcell_out_25[2] dcim_bitcell
xi_bitcell_25_3 vdd gnd wl[25] in_b[25] bl[3] bl_b[3] bitcell_out_25[3] dcim_bitcell
xi_bitcell_26_0 vdd gnd wl[26] in_b[26] bl[0] bl_b[0] bitcell_out_26[0] dcim_bitcell
xi_bitcell_26_1 vdd gnd wl[26] in_b[26] bl[1] bl_b[1] bitcell_out_26[1] dcim_bitcell
xi_bitcell_26_2 vdd gnd wl[26] in_b[26] bl[2] bl_b[2] bitcell_out_26[2] dcim_bitcell
xi_bitcell_26_3 vdd gnd wl[26] in_b[26] bl[3] bl_b[3] bitcell_out_26[3] dcim_bitcell
xi_bitcell_27_0 vdd gnd wl[27] in_b[27] bl[0] bl_b[0] bitcell_out_27[0] dcim_bitcell
xi_bitcell_27_1 vdd gnd wl[27] in_b[27] bl[1] bl_b[1] bitcell_out_27[1] dcim_bitcell
xi_bitcell_27_2 vdd gnd wl[27] in_b[27] bl[2] bl_b[2] bitcell_out_27[2] dcim_bitcell
xi_bitcell_27_3 vdd gnd wl[27] in_b[27] bl[3] bl_b[3] bitcell_out_27[3] dcim_bitcell
xi_bitcell_28_0 vdd gnd wl[28] in_b[28] bl[0] bl_b[0] bitcell_out_28[0] dcim_bitcell
xi_bitcell_28_1 vdd gnd wl[28] in_b[28] bl[1] bl_b[1] bitcell_out_28[1] dcim_bitcell
xi_bitcell_28_2 vdd gnd wl[28] in_b[28] bl[2] bl_b[2] bitcell_out_28[2] dcim_bitcell
xi_bitcell_28_3 vdd gnd wl[28] in_b[28] bl[3] bl_b[3] bitcell_out_28[3] dcim_bitcell
xi_bitcell_29_0 vdd gnd wl[29] in_b[29] bl[0] bl_b[0] bitcell_out_29[0] dcim_bitcell
xi_bitcell_29_1 vdd gnd wl[29] in_b[29] bl[1] bl_b[1] bitcell_out_29[1] dcim_bitcell
xi_bitcell_29_2 vdd gnd wl[29] in_b[29] bl[2] bl_b[2] bitcell_out_29[2] dcim_bitcell
xi_bitcell_29_3 vdd gnd wl[29] in_b[29] bl[3] bl_b[3] bitcell_out_29[3] dcim_bitcell
xi_bitcell_30_0 vdd gnd wl[30] in_b[30] bl[0] bl_b[0] bitcell_out_30[0] dcim_bitcell
xi_bitcell_30_1 vdd gnd wl[30] in_b[30] bl[1] bl_b[1] bitcell_out_30[1] dcim_bitcell
xi_bitcell_30_2 vdd gnd wl[30] in_b[30] bl[2] bl_b[2] bitcell_out_30[2] dcim_bitcell
xi_bitcell_30_3 vdd gnd wl[30] in_b[30] bl[3] bl_b[3] bitcell_out_30[3] dcim_bitcell
xi_bitcell_31_0 vdd gnd wl[31] in_b[31] bl[0] bl_b[0] bitcell_out_31[0] dcim_bitcell
xi_bitcell_31_1 vdd gnd wl[31] in_b[31] bl[1] bl_b[1] bitcell_out_31[1] dcim_bitcell
xi_bitcell_31_2 vdd gnd wl[31] in_b[31] bl[2] bl_b[2] bitcell_out_31[2] dcim_bitcell
xi_bitcell_31_3 vdd gnd wl[31] in_b[31] bl[3] bl_b[3] bitcell_out_31[3] dcim_bitcell
xi_bitcell_32_0 vdd gnd wl[32] in_b[32] bl[0] bl_b[0] bitcell_out_32[0] dcim_bitcell
xi_bitcell_32_1 vdd gnd wl[32] in_b[32] bl[1] bl_b[1] bitcell_out_32[1] dcim_bitcell
xi_bitcell_32_2 vdd gnd wl[32] in_b[32] bl[2] bl_b[2] bitcell_out_32[2] dcim_bitcell
xi_bitcell_32_3 vdd gnd wl[32] in_b[32] bl[3] bl_b[3] bitcell_out_32[3] dcim_bitcell
xi_bitcell_33_0 vdd gnd wl[33] in_b[33] bl[0] bl_b[0] bitcell_out_33[0] dcim_bitcell
xi_bitcell_33_1 vdd gnd wl[33] in_b[33] bl[1] bl_b[1] bitcell_out_33[1] dcim_bitcell
xi_bitcell_33_2 vdd gnd wl[33] in_b[33] bl[2] bl_b[2] bitcell_out_33[2] dcim_bitcell
xi_bitcell_33_3 vdd gnd wl[33] in_b[33] bl[3] bl_b[3] bitcell_out_33[3] dcim_bitcell
xi_bitcell_34_0 vdd gnd wl[34] in_b[34] bl[0] bl_b[0] bitcell_out_34[0] dcim_bitcell
xi_bitcell_34_1 vdd gnd wl[34] in_b[34] bl[1] bl_b[1] bitcell_out_34[1] dcim_bitcell
xi_bitcell_34_2 vdd gnd wl[34] in_b[34] bl[2] bl_b[2] bitcell_out_34[2] dcim_bitcell
xi_bitcell_34_3 vdd gnd wl[34] in_b[34] bl[3] bl_b[3] bitcell_out_34[3] dcim_bitcell
xi_bitcell_35_0 vdd gnd wl[35] in_b[35] bl[0] bl_b[0] bitcell_out_35[0] dcim_bitcell
xi_bitcell_35_1 vdd gnd wl[35] in_b[35] bl[1] bl_b[1] bitcell_out_35[1] dcim_bitcell
xi_bitcell_35_2 vdd gnd wl[35] in_b[35] bl[2] bl_b[2] bitcell_out_35[2] dcim_bitcell
xi_bitcell_35_3 vdd gnd wl[35] in_b[35] bl[3] bl_b[3] bitcell_out_35[3] dcim_bitcell
xi_bitcell_36_0 vdd gnd wl[36] in_b[36] bl[0] bl_b[0] bitcell_out_36[0] dcim_bitcell
xi_bitcell_36_1 vdd gnd wl[36] in_b[36] bl[1] bl_b[1] bitcell_out_36[1] dcim_bitcell
xi_bitcell_36_2 vdd gnd wl[36] in_b[36] bl[2] bl_b[2] bitcell_out_36[2] dcim_bitcell
xi_bitcell_36_3 vdd gnd wl[36] in_b[36] bl[3] bl_b[3] bitcell_out_36[3] dcim_bitcell
xi_bitcell_37_0 vdd gnd wl[37] in_b[37] bl[0] bl_b[0] bitcell_out_37[0] dcim_bitcell
xi_bitcell_37_1 vdd gnd wl[37] in_b[37] bl[1] bl_b[1] bitcell_out_37[1] dcim_bitcell
xi_bitcell_37_2 vdd gnd wl[37] in_b[37] bl[2] bl_b[2] bitcell_out_37[2] dcim_bitcell
xi_bitcell_37_3 vdd gnd wl[37] in_b[37] bl[3] bl_b[3] bitcell_out_37[3] dcim_bitcell
xi_bitcell_38_0 vdd gnd wl[38] in_b[38] bl[0] bl_b[0] bitcell_out_38[0] dcim_bitcell
xi_bitcell_38_1 vdd gnd wl[38] in_b[38] bl[1] bl_b[1] bitcell_out_38[1] dcim_bitcell
xi_bitcell_38_2 vdd gnd wl[38] in_b[38] bl[2] bl_b[2] bitcell_out_38[2] dcim_bitcell
xi_bitcell_38_3 vdd gnd wl[38] in_b[38] bl[3] bl_b[3] bitcell_out_38[3] dcim_bitcell
xi_bitcell_39_0 vdd gnd wl[39] in_b[39] bl[0] bl_b[0] bitcell_out_39[0] dcim_bitcell
xi_bitcell_39_1 vdd gnd wl[39] in_b[39] bl[1] bl_b[1] bitcell_out_39[1] dcim_bitcell
xi_bitcell_39_2 vdd gnd wl[39] in_b[39] bl[2] bl_b[2] bitcell_out_39[2] dcim_bitcell
xi_bitcell_39_3 vdd gnd wl[39] in_b[39] bl[3] bl_b[3] bitcell_out_39[3] dcim_bitcell
xi_bitcell_40_0 vdd gnd wl[40] in_b[40] bl[0] bl_b[0] bitcell_out_40[0] dcim_bitcell
xi_bitcell_40_1 vdd gnd wl[40] in_b[40] bl[1] bl_b[1] bitcell_out_40[1] dcim_bitcell
xi_bitcell_40_2 vdd gnd wl[40] in_b[40] bl[2] bl_b[2] bitcell_out_40[2] dcim_bitcell
xi_bitcell_40_3 vdd gnd wl[40] in_b[40] bl[3] bl_b[3] bitcell_out_40[3] dcim_bitcell
xi_bitcell_41_0 vdd gnd wl[41] in_b[41] bl[0] bl_b[0] bitcell_out_41[0] dcim_bitcell
xi_bitcell_41_1 vdd gnd wl[41] in_b[41] bl[1] bl_b[1] bitcell_out_41[1] dcim_bitcell
xi_bitcell_41_2 vdd gnd wl[41] in_b[41] bl[2] bl_b[2] bitcell_out_41[2] dcim_bitcell
xi_bitcell_41_3 vdd gnd wl[41] in_b[41] bl[3] bl_b[3] bitcell_out_41[3] dcim_bitcell
xi_bitcell_42_0 vdd gnd wl[42] in_b[42] bl[0] bl_b[0] bitcell_out_42[0] dcim_bitcell
xi_bitcell_42_1 vdd gnd wl[42] in_b[42] bl[1] bl_b[1] bitcell_out_42[1] dcim_bitcell
xi_bitcell_42_2 vdd gnd wl[42] in_b[42] bl[2] bl_b[2] bitcell_out_42[2] dcim_bitcell
xi_bitcell_42_3 vdd gnd wl[42] in_b[42] bl[3] bl_b[3] bitcell_out_42[3] dcim_bitcell
xi_bitcell_43_0 vdd gnd wl[43] in_b[43] bl[0] bl_b[0] bitcell_out_43[0] dcim_bitcell
xi_bitcell_43_1 vdd gnd wl[43] in_b[43] bl[1] bl_b[1] bitcell_out_43[1] dcim_bitcell
xi_bitcell_43_2 vdd gnd wl[43] in_b[43] bl[2] bl_b[2] bitcell_out_43[2] dcim_bitcell
xi_bitcell_43_3 vdd gnd wl[43] in_b[43] bl[3] bl_b[3] bitcell_out_43[3] dcim_bitcell
xi_bitcell_44_0 vdd gnd wl[44] in_b[44] bl[0] bl_b[0] bitcell_out_44[0] dcim_bitcell
xi_bitcell_44_1 vdd gnd wl[44] in_b[44] bl[1] bl_b[1] bitcell_out_44[1] dcim_bitcell
xi_bitcell_44_2 vdd gnd wl[44] in_b[44] bl[2] bl_b[2] bitcell_out_44[2] dcim_bitcell
xi_bitcell_44_3 vdd gnd wl[44] in_b[44] bl[3] bl_b[3] bitcell_out_44[3] dcim_bitcell
xi_bitcell_45_0 vdd gnd wl[45] in_b[45] bl[0] bl_b[0] bitcell_out_45[0] dcim_bitcell
xi_bitcell_45_1 vdd gnd wl[45] in_b[45] bl[1] bl_b[1] bitcell_out_45[1] dcim_bitcell
xi_bitcell_45_2 vdd gnd wl[45] in_b[45] bl[2] bl_b[2] bitcell_out_45[2] dcim_bitcell
xi_bitcell_45_3 vdd gnd wl[45] in_b[45] bl[3] bl_b[3] bitcell_out_45[3] dcim_bitcell
xi_bitcell_46_0 vdd gnd wl[46] in_b[46] bl[0] bl_b[0] bitcell_out_46[0] dcim_bitcell
xi_bitcell_46_1 vdd gnd wl[46] in_b[46] bl[1] bl_b[1] bitcell_out_46[1] dcim_bitcell
xi_bitcell_46_2 vdd gnd wl[46] in_b[46] bl[2] bl_b[2] bitcell_out_46[2] dcim_bitcell
xi_bitcell_46_3 vdd gnd wl[46] in_b[46] bl[3] bl_b[3] bitcell_out_46[3] dcim_bitcell
xi_bitcell_47_0 vdd gnd wl[47] in_b[47] bl[0] bl_b[0] bitcell_out_47[0] dcim_bitcell
xi_bitcell_47_1 vdd gnd wl[47] in_b[47] bl[1] bl_b[1] bitcell_out_47[1] dcim_bitcell
xi_bitcell_47_2 vdd gnd wl[47] in_b[47] bl[2] bl_b[2] bitcell_out_47[2] dcim_bitcell
xi_bitcell_47_3 vdd gnd wl[47] in_b[47] bl[3] bl_b[3] bitcell_out_47[3] dcim_bitcell
xi_bitcell_48_0 vdd gnd wl[48] in_b[48] bl[0] bl_b[0] bitcell_out_48[0] dcim_bitcell
xi_bitcell_48_1 vdd gnd wl[48] in_b[48] bl[1] bl_b[1] bitcell_out_48[1] dcim_bitcell
xi_bitcell_48_2 vdd gnd wl[48] in_b[48] bl[2] bl_b[2] bitcell_out_48[2] dcim_bitcell
xi_bitcell_48_3 vdd gnd wl[48] in_b[48] bl[3] bl_b[3] bitcell_out_48[3] dcim_bitcell
xi_bitcell_49_0 vdd gnd wl[49] in_b[49] bl[0] bl_b[0] bitcell_out_49[0] dcim_bitcell
xi_bitcell_49_1 vdd gnd wl[49] in_b[49] bl[1] bl_b[1] bitcell_out_49[1] dcim_bitcell
xi_bitcell_49_2 vdd gnd wl[49] in_b[49] bl[2] bl_b[2] bitcell_out_49[2] dcim_bitcell
xi_bitcell_49_3 vdd gnd wl[49] in_b[49] bl[3] bl_b[3] bitcell_out_49[3] dcim_bitcell
xi_bitcell_50_0 vdd gnd wl[50] in_b[50] bl[0] bl_b[0] bitcell_out_50[0] dcim_bitcell
xi_bitcell_50_1 vdd gnd wl[50] in_b[50] bl[1] bl_b[1] bitcell_out_50[1] dcim_bitcell
xi_bitcell_50_2 vdd gnd wl[50] in_b[50] bl[2] bl_b[2] bitcell_out_50[2] dcim_bitcell
xi_bitcell_50_3 vdd gnd wl[50] in_b[50] bl[3] bl_b[3] bitcell_out_50[3] dcim_bitcell
xi_bitcell_51_0 vdd gnd wl[51] in_b[51] bl[0] bl_b[0] bitcell_out_51[0] dcim_bitcell
xi_bitcell_51_1 vdd gnd wl[51] in_b[51] bl[1] bl_b[1] bitcell_out_51[1] dcim_bitcell
xi_bitcell_51_2 vdd gnd wl[51] in_b[51] bl[2] bl_b[2] bitcell_out_51[2] dcim_bitcell
xi_bitcell_51_3 vdd gnd wl[51] in_b[51] bl[3] bl_b[3] bitcell_out_51[3] dcim_bitcell
xi_bitcell_52_0 vdd gnd wl[52] in_b[52] bl[0] bl_b[0] bitcell_out_52[0] dcim_bitcell
xi_bitcell_52_1 vdd gnd wl[52] in_b[52] bl[1] bl_b[1] bitcell_out_52[1] dcim_bitcell
xi_bitcell_52_2 vdd gnd wl[52] in_b[52] bl[2] bl_b[2] bitcell_out_52[2] dcim_bitcell
xi_bitcell_52_3 vdd gnd wl[52] in_b[52] bl[3] bl_b[3] bitcell_out_52[3] dcim_bitcell
xi_bitcell_53_0 vdd gnd wl[53] in_b[53] bl[0] bl_b[0] bitcell_out_53[0] dcim_bitcell
xi_bitcell_53_1 vdd gnd wl[53] in_b[53] bl[1] bl_b[1] bitcell_out_53[1] dcim_bitcell
xi_bitcell_53_2 vdd gnd wl[53] in_b[53] bl[2] bl_b[2] bitcell_out_53[2] dcim_bitcell
xi_bitcell_53_3 vdd gnd wl[53] in_b[53] bl[3] bl_b[3] bitcell_out_53[3] dcim_bitcell
xi_bitcell_54_0 vdd gnd wl[54] in_b[54] bl[0] bl_b[0] bitcell_out_54[0] dcim_bitcell
xi_bitcell_54_1 vdd gnd wl[54] in_b[54] bl[1] bl_b[1] bitcell_out_54[1] dcim_bitcell
xi_bitcell_54_2 vdd gnd wl[54] in_b[54] bl[2] bl_b[2] bitcell_out_54[2] dcim_bitcell
xi_bitcell_54_3 vdd gnd wl[54] in_b[54] bl[3] bl_b[3] bitcell_out_54[3] dcim_bitcell
xi_bitcell_55_0 vdd gnd wl[55] in_b[55] bl[0] bl_b[0] bitcell_out_55[0] dcim_bitcell
xi_bitcell_55_1 vdd gnd wl[55] in_b[55] bl[1] bl_b[1] bitcell_out_55[1] dcim_bitcell
xi_bitcell_55_2 vdd gnd wl[55] in_b[55] bl[2] bl_b[2] bitcell_out_55[2] dcim_bitcell
xi_bitcell_55_3 vdd gnd wl[55] in_b[55] bl[3] bl_b[3] bitcell_out_55[3] dcim_bitcell
xi_bitcell_56_0 vdd gnd wl[56] in_b[56] bl[0] bl_b[0] bitcell_out_56[0] dcim_bitcell
xi_bitcell_56_1 vdd gnd wl[56] in_b[56] bl[1] bl_b[1] bitcell_out_56[1] dcim_bitcell
xi_bitcell_56_2 vdd gnd wl[56] in_b[56] bl[2] bl_b[2] bitcell_out_56[2] dcim_bitcell
xi_bitcell_56_3 vdd gnd wl[56] in_b[56] bl[3] bl_b[3] bitcell_out_56[3] dcim_bitcell
xi_bitcell_57_0 vdd gnd wl[57] in_b[57] bl[0] bl_b[0] bitcell_out_57[0] dcim_bitcell
xi_bitcell_57_1 vdd gnd wl[57] in_b[57] bl[1] bl_b[1] bitcell_out_57[1] dcim_bitcell
xi_bitcell_57_2 vdd gnd wl[57] in_b[57] bl[2] bl_b[2] bitcell_out_57[2] dcim_bitcell
xi_bitcell_57_3 vdd gnd wl[57] in_b[57] bl[3] bl_b[3] bitcell_out_57[3] dcim_bitcell
xi_bitcell_58_0 vdd gnd wl[58] in_b[58] bl[0] bl_b[0] bitcell_out_58[0] dcim_bitcell
xi_bitcell_58_1 vdd gnd wl[58] in_b[58] bl[1] bl_b[1] bitcell_out_58[1] dcim_bitcell
xi_bitcell_58_2 vdd gnd wl[58] in_b[58] bl[2] bl_b[2] bitcell_out_58[2] dcim_bitcell
xi_bitcell_58_3 vdd gnd wl[58] in_b[58] bl[3] bl_b[3] bitcell_out_58[3] dcim_bitcell
xi_bitcell_59_0 vdd gnd wl[59] in_b[59] bl[0] bl_b[0] bitcell_out_59[0] dcim_bitcell
xi_bitcell_59_1 vdd gnd wl[59] in_b[59] bl[1] bl_b[1] bitcell_out_59[1] dcim_bitcell
xi_bitcell_59_2 vdd gnd wl[59] in_b[59] bl[2] bl_b[2] bitcell_out_59[2] dcim_bitcell
xi_bitcell_59_3 vdd gnd wl[59] in_b[59] bl[3] bl_b[3] bitcell_out_59[3] dcim_bitcell
xi_bitcell_60_0 vdd gnd wl[60] in_b[60] bl[0] bl_b[0] bitcell_out_60[0] dcim_bitcell
xi_bitcell_60_1 vdd gnd wl[60] in_b[60] bl[1] bl_b[1] bitcell_out_60[1] dcim_bitcell
xi_bitcell_60_2 vdd gnd wl[60] in_b[60] bl[2] bl_b[2] bitcell_out_60[2] dcim_bitcell
xi_bitcell_60_3 vdd gnd wl[60] in_b[60] bl[3] bl_b[3] bitcell_out_60[3] dcim_bitcell
xi_bitcell_61_0 vdd gnd wl[61] in_b[61] bl[0] bl_b[0] bitcell_out_61[0] dcim_bitcell
xi_bitcell_61_1 vdd gnd wl[61] in_b[61] bl[1] bl_b[1] bitcell_out_61[1] dcim_bitcell
xi_bitcell_61_2 vdd gnd wl[61] in_b[61] bl[2] bl_b[2] bitcell_out_61[2] dcim_bitcell
xi_bitcell_61_3 vdd gnd wl[61] in_b[61] bl[3] bl_b[3] bitcell_out_61[3] dcim_bitcell
xi_bitcell_62_0 vdd gnd wl[62] in_b[62] bl[0] bl_b[0] bitcell_out_62[0] dcim_bitcell
xi_bitcell_62_1 vdd gnd wl[62] in_b[62] bl[1] bl_b[1] bitcell_out_62[1] dcim_bitcell
xi_bitcell_62_2 vdd gnd wl[62] in_b[62] bl[2] bl_b[2] bitcell_out_62[2] dcim_bitcell
xi_bitcell_62_3 vdd gnd wl[62] in_b[62] bl[3] bl_b[3] bitcell_out_62[3] dcim_bitcell
xi_bitcell_63_0 vdd gnd wl[63] in_b[63] bl[0] bl_b[0] bitcell_out_63[0] dcim_bitcell
xi_bitcell_63_1 vdd gnd wl[63] in_b[63] bl[1] bl_b[1] bitcell_out_63[1] dcim_bitcell
xi_bitcell_63_2 vdd gnd wl[63] in_b[63] bl[2] bl_b[2] bitcell_out_63[2] dcim_bitcell
xi_bitcell_63_3 vdd gnd wl[63] in_b[63] bl[3] bl_b[3] bitcell_out_63[3] dcim_bitcell
.ends sram_64x4
** End of subcircuit definition.

** Cell name: sram_rw_4bit
.subckt sram_rw_4bit vdd gnd bl[0] bl[1] bl[2] bl[3] bl_b[0] bl_b[1] bl_b[2] bl_b[3] pe ysw ysr spe se din[0] din[1] din[2] din[3] dout[0] dout[1] dout[2] dout[3] 
xi_rw_0 vdd gnd bl[0] bl_b[0] pe ysw ysr spe se din[0] dout[0] sram_rw
xi_rw_1 vdd gnd bl[1] bl_b[1] pe ysw ysr spe se din[1] dout[1] sram_rw
xi_rw_2 vdd gnd bl[2] bl_b[2] pe ysw ysr spe se din[2] dout[2] sram_rw
xi_rw_3 vdd gnd bl[3] bl_b[3] pe ysw ysr spe se din[3] dout[3] sram_rw
.ends sram_rw_4bit
** End of subcircuit definition.

** Cell name: sram_64x4_with_rw
.subckt sram_64x4_with_rw vdd gnd pe ysw ysr spe se wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] in_b[0] in_b[1] in_b[2] in_b[3] in_b[4] in_b[5] in_b[6] in_b[7] in_b[8] in_b[9] in_b[10] in_b[11] in_b[12] in_b[13] in_b[14] in_b[15] in_b[16] in_b[17] in_b[18] in_b[19] in_b[20] in_b[21] in_b[22] in_b[23] in_b[24] in_b[25] in_b[26] in_b[27] in_b[28] in_b[29] in_b[30] in_b[31] in_b[32] in_b[33] in_b[34] in_b[35] in_b[36] in_b[37] in_b[38] in_b[39] in_b[40] in_b[41] in_b[42] in_b[43] in_b[44] in_b[45] in_b[46] in_b[47] in_b[48] in_b[49] in_b[50] in_b[51] in_b[52] in_b[53] in_b[54] in_b[55] in_b[56] in_b[57] in_b[58] in_b[59] in_b[60] in_b[61] in_b[62] in_b[63] din[0] din[1] din[2] din[3] dout[0] dout[1] dout[2] dout[3] bitcell_out_0[0] bitcell_out_0[1] bitcell_out_0[2] bitcell_out_0[3] bitcell_out_1[0] bitcell_out_1[1] bitcell_out_1[2] bitcell_out_1[3] bitcell_out_2[0] bitcell_out_2[1] bitcell_out_2[2] bitcell_out_2[3] bitcell_out_3[0] bitcell_out_3[1] bitcell_out_3[2] bitcell_out_3[3] bitcell_out_4[0] bitcell_out_4[1] bitcell_out_4[2] bitcell_out_4[3] bitcell_out_5[0] bitcell_out_5[1] bitcell_out_5[2] bitcell_out_5[3] bitcell_out_6[0] bitcell_out_6[1] bitcell_out_6[2] bitcell_out_6[3] bitcell_out_7[0] bitcell_out_7[1] bitcell_out_7[2] bitcell_out_7[3] bitcell_out_8[0] bitcell_out_8[1] bitcell_out_8[2] bitcell_out_8[3] bitcell_out_9[0] bitcell_out_9[1] bitcell_out_9[2] bitcell_out_9[3] bitcell_out_10[0] bitcell_out_10[1] bitcell_out_10[2] bitcell_out_10[3] bitcell_out_11[0] bitcell_out_11[1] bitcell_out_11[2] bitcell_out_11[3] bitcell_out_12[0] bitcell_out_12[1] bitcell_out_12[2] bitcell_out_12[3] bitcell_out_13[0] bitcell_out_13[1] bitcell_out_13[2] bitcell_out_13[3] bitcell_out_14[0] bitcell_out_14[1] bitcell_out_14[2] bitcell_out_14[3] bitcell_out_15[0] bitcell_out_15[1] bitcell_out_15[2] bitcell_out_15[3] bitcell_out_16[0] bitcell_out_16[1] bitcell_out_16[2] bitcell_out_16[3] bitcell_out_17[0] bitcell_out_17[1] bitcell_out_17[2] bitcell_out_17[3] bitcell_out_18[0] bitcell_out_18[1] bitcell_out_18[2] bitcell_out_18[3] bitcell_out_19[0] bitcell_out_19[1] bitcell_out_19[2] bitcell_out_19[3] bitcell_out_20[0] bitcell_out_20[1] bitcell_out_20[2] bitcell_out_20[3] bitcell_out_21[0] bitcell_out_21[1] bitcell_out_21[2] bitcell_out_21[3] bitcell_out_22[0] bitcell_out_22[1] bitcell_out_22[2] bitcell_out_22[3] bitcell_out_23[0] bitcell_out_23[1] bitcell_out_23[2] bitcell_out_23[3] bitcell_out_24[0] bitcell_out_24[1] bitcell_out_24[2] bitcell_out_24[3] bitcell_out_25[0] bitcell_out_25[1] bitcell_out_25[2] bitcell_out_25[3] bitcell_out_26[0] bitcell_out_26[1] bitcell_out_26[2] bitcell_out_26[3] bitcell_out_27[0] bitcell_out_27[1] bitcell_out_27[2] bitcell_out_27[3] bitcell_out_28[0] bitcell_out_28[1] bitcell_out_28[2] bitcell_out_28[3] bitcell_out_29[0] bitcell_out_29[1] bitcell_out_29[2] bitcell_out_29[3] bitcell_out_30[0] bitcell_out_30[1] bitcell_out_30[2] bitcell_out_30[3] bitcell_out_31[0] bitcell_out_31[1] bitcell_out_31[2] bitcell_out_31[3] bitcell_out_32[0] bitcell_out_32[1] bitcell_out_32[2] bitcell_out_32[3] bitcell_out_33[0] bitcell_out_33[1] bitcell_out_33[2] bitcell_out_33[3] bitcell_out_34[0] bitcell_out_34[1] bitcell_out_34[2] bitcell_out_34[3] bitcell_out_35[0] bitcell_out_35[1] bitcell_out_35[2] bitcell_out_35[3] bitcell_out_36[0] bitcell_out_36[1] bitcell_out_36[2] bitcell_out_36[3] bitcell_out_37[0] bitcell_out_37[1] bitcell_out_37[2] bitcell_out_37[3] bitcell_out_38[0] bitcell_out_38[1] bitcell_out_38[2] bitcell_out_38[3] bitcell_out_39[0] bitcell_out_39[1] bitcell_out_39[2] bitcell_out_39[3] bitcell_out_40[0] bitcell_out_40[1] bitcell_out_40[2] bitcell_out_40[3] bitcell_out_41[0] bitcell_out_41[1] bitcell_out_41[2] bitcell_out_41[3] bitcell_out_42[0] bitcell_out_42[1] bitcell_out_42[2] bitcell_out_42[3] bitcell_out_43[0] bitcell_out_43[1] bitcell_out_43[2] bitcell_out_43[3] bitcell_out_44[0] bitcell_out_44[1] bitcell_out_44[2] bitcell_out_44[3] bitcell_out_45[0] bitcell_out_45[1] bitcell_out_45[2] bitcell_out_45[3] bitcell_out_46[0] bitcell_out_46[1] bitcell_out_46[2] bitcell_out_46[3] bitcell_out_47[0] bitcell_out_47[1] bitcell_out_47[2] bitcell_out_47[3] bitcell_out_48[0] bitcell_out_48[1] bitcell_out_48[2] bitcell_out_48[3] bitcell_out_49[0] bitcell_out_49[1] bitcell_out_49[2] bitcell_out_49[3] bitcell_out_50[0] bitcell_out_50[1] bitcell_out_50[2] bitcell_out_50[3] bitcell_out_51[0] bitcell_out_51[1] bitcell_out_51[2] bitcell_out_51[3] bitcell_out_52[0] bitcell_out_52[1] bitcell_out_52[2] bitcell_out_52[3] bitcell_out_53[0] bitcell_out_53[1] bitcell_out_53[2] bitcell_out_53[3] bitcell_out_54[0] bitcell_out_54[1] bitcell_out_54[2] bitcell_out_54[3] bitcell_out_55[0] bitcell_out_55[1] bitcell_out_55[2] bitcell_out_55[3] bitcell_out_56[0] bitcell_out_56[1] bitcell_out_56[2] bitcell_out_56[3] bitcell_out_57[0] bitcell_out_57[1] bitcell_out_57[2] bitcell_out_57[3] bitcell_out_58[0] bitcell_out_58[1] bitcell_out_58[2] bitcell_out_58[3] bitcell_out_59[0] bitcell_out_59[1] bitcell_out_59[2] bitcell_out_59[3] bitcell_out_60[0] bitcell_out_60[1] bitcell_out_60[2] bitcell_out_60[3] bitcell_out_61[0] bitcell_out_61[1] bitcell_out_61[2] bitcell_out_61[3] bitcell_out_62[0] bitcell_out_62[1] bitcell_out_62[2] bitcell_out_62[3] bitcell_out_63[0] bitcell_out_63[1] bitcell_out_63[2] bitcell_out_63[3] 
xi_sram vdd gnd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] in_b[0] in_b[1] in_b[2] in_b[3] in_b[4] in_b[5] in_b[6] in_b[7] in_b[8] in_b[9] in_b[10] in_b[11] in_b[12] in_b[13] in_b[14] in_b[15] in_b[16] in_b[17] in_b[18] in_b[19] in_b[20] in_b[21] in_b[22] in_b[23] in_b[24] in_b[25] in_b[26] in_b[27] in_b[28] in_b[29] in_b[30] in_b[31] in_b[32] in_b[33] in_b[34] in_b[35] in_b[36] in_b[37] in_b[38] in_b[39] in_b[40] in_b[41] in_b[42] in_b[43] in_b[44] in_b[45] in_b[46] in_b[47] in_b[48] in_b[49] in_b[50] in_b[51] in_b[52] in_b[53] in_b[54] in_b[55] in_b[56] in_b[57] in_b[58] in_b[59] in_b[60] in_b[61] in_b[62] in_b[63] bl[0] bl[1] bl[2] bl[3] bl_b[0] bl_b[1] bl_b[2] bl_b[3] bitcell_out_0[0] bitcell_out_0[1] bitcell_out_0[2] bitcell_out_0[3] bitcell_out_1[0] bitcell_out_1[1] bitcell_out_1[2] bitcell_out_1[3] bitcell_out_2[0] bitcell_out_2[1] bitcell_out_2[2] bitcell_out_2[3] bitcell_out_3[0] bitcell_out_3[1] bitcell_out_3[2] bitcell_out_3[3] bitcell_out_4[0] bitcell_out_4[1] bitcell_out_4[2] bitcell_out_4[3] bitcell_out_5[0] bitcell_out_5[1] bitcell_out_5[2] bitcell_out_5[3] bitcell_out_6[0] bitcell_out_6[1] bitcell_out_6[2] bitcell_out_6[3] bitcell_out_7[0] bitcell_out_7[1] bitcell_out_7[2] bitcell_out_7[3] bitcell_out_8[0] bitcell_out_8[1] bitcell_out_8[2] bitcell_out_8[3] bitcell_out_9[0] bitcell_out_9[1] bitcell_out_9[2] bitcell_out_9[3] bitcell_out_10[0] bitcell_out_10[1] bitcell_out_10[2] bitcell_out_10[3] bitcell_out_11[0] bitcell_out_11[1] bitcell_out_11[2] bitcell_out_11[3] bitcell_out_12[0] bitcell_out_12[1] bitcell_out_12[2] bitcell_out_12[3] bitcell_out_13[0] bitcell_out_13[1] bitcell_out_13[2] bitcell_out_13[3] bitcell_out_14[0] bitcell_out_14[1] bitcell_out_14[2] bitcell_out_14[3] bitcell_out_15[0] bitcell_out_15[1] bitcell_out_15[2] bitcell_out_15[3] bitcell_out_16[0] bitcell_out_16[1] bitcell_out_16[2] bitcell_out_16[3] bitcell_out_17[0] bitcell_out_17[1] bitcell_out_17[2] bitcell_out_17[3] bitcell_out_18[0] bitcell_out_18[1] bitcell_out_18[2] bitcell_out_18[3] bitcell_out_19[0] bitcell_out_19[1] bitcell_out_19[2] bitcell_out_19[3] bitcell_out_20[0] bitcell_out_20[1] bitcell_out_20[2] bitcell_out_20[3] bitcell_out_21[0] bitcell_out_21[1] bitcell_out_21[2] bitcell_out_21[3] bitcell_out_22[0] bitcell_out_22[1] bitcell_out_22[2] bitcell_out_22[3] bitcell_out_23[0] bitcell_out_23[1] bitcell_out_23[2] bitcell_out_23[3] bitcell_out_24[0] bitcell_out_24[1] bitcell_out_24[2] bitcell_out_24[3] bitcell_out_25[0] bitcell_out_25[1] bitcell_out_25[2] bitcell_out_25[3] bitcell_out_26[0] bitcell_out_26[1] bitcell_out_26[2] bitcell_out_26[3] bitcell_out_27[0] bitcell_out_27[1] bitcell_out_27[2] bitcell_out_27[3] bitcell_out_28[0] bitcell_out_28[1] bitcell_out_28[2] bitcell_out_28[3] bitcell_out_29[0] bitcell_out_29[1] bitcell_out_29[2] bitcell_out_29[3] bitcell_out_30[0] bitcell_out_30[1] bitcell_out_30[2] bitcell_out_30[3] bitcell_out_31[0] bitcell_out_31[1] bitcell_out_31[2] bitcell_out_31[3] bitcell_out_32[0] bitcell_out_32[1] bitcell_out_32[2] bitcell_out_32[3] bitcell_out_33[0] bitcell_out_33[1] bitcell_out_33[2] bitcell_out_33[3] bitcell_out_34[0] bitcell_out_34[1] bitcell_out_34[2] bitcell_out_34[3] bitcell_out_35[0] bitcell_out_35[1] bitcell_out_35[2] bitcell_out_35[3] bitcell_out_36[0] bitcell_out_36[1] bitcell_out_36[2] bitcell_out_36[3] bitcell_out_37[0] bitcell_out_37[1] bitcell_out_37[2] bitcell_out_37[3] bitcell_out_38[0] bitcell_out_38[1] bitcell_out_38[2] bitcell_out_38[3] bitcell_out_39[0] bitcell_out_39[1] bitcell_out_39[2] bitcell_out_39[3] bitcell_out_40[0] bitcell_out_40[1] bitcell_out_40[2] bitcell_out_40[3] bitcell_out_41[0] bitcell_out_41[1] bitcell_out_41[2] bitcell_out_41[3] bitcell_out_42[0] bitcell_out_42[1] bitcell_out_42[2] bitcell_out_42[3] bitcell_out_43[0] bitcell_out_43[1] bitcell_out_43[2] bitcell_out_43[3] bitcell_out_44[0] bitcell_out_44[1] bitcell_out_44[2] bitcell_out_44[3] bitcell_out_45[0] bitcell_out_45[1] bitcell_out_45[2] bitcell_out_45[3] bitcell_out_46[0] bitcell_out_46[1] bitcell_out_46[2] bitcell_out_46[3] bitcell_out_47[0] bitcell_out_47[1] bitcell_out_47[2] bitcell_out_47[3] bitcell_out_48[0] bitcell_out_48[1] bitcell_out_48[2] bitcell_out_48[3] bitcell_out_49[0] bitcell_out_49[1] bitcell_out_49[2] bitcell_out_49[3] bitcell_out_50[0] bitcell_out_50[1] bitcell_out_50[2] bitcell_out_50[3] bitcell_out_51[0] bitcell_out_51[1] bitcell_out_51[2] bitcell_out_51[3] bitcell_out_52[0] bitcell_out_52[1] bitcell_out_52[2] bitcell_out_52[3] bitcell_out_53[0] bitcell_out_53[1] bitcell_out_53[2] bitcell_out_53[3] bitcell_out_54[0] bitcell_out_54[1] bitcell_out_54[2] bitcell_out_54[3] bitcell_out_55[0] bitcell_out_55[1] bitcell_out_55[2] bitcell_out_55[3] bitcell_out_56[0] bitcell_out_56[1] bitcell_out_56[2] bitcell_out_56[3] bitcell_out_57[0] bitcell_out_57[1] bitcell_out_57[2] bitcell_out_57[3] bitcell_out_58[0] bitcell_out_58[1] bitcell_out_58[2] bitcell_out_58[3] bitcell_out_59[0] bitcell_out_59[1] bitcell_out_59[2] bitcell_out_59[3] bitcell_out_60[0] bitcell_out_60[1] bitcell_out_60[2] bitcell_out_60[3] bitcell_out_61[0] bitcell_out_61[1] bitcell_out_61[2] bitcell_out_61[3] bitcell_out_62[0] bitcell_out_62[1] bitcell_out_62[2] bitcell_out_62[3] bitcell_out_63[0] bitcell_out_63[1] bitcell_out_63[2] bitcell_out_63[3] sram_64x4
xi_sram_rw vdd gnd bl[0] bl[1] bl[2] bl[3] bl_b[0] bl_b[1] bl_b[2] bl_b[3] pe ysw ysr spe se din[0] din[1] din[2] din[3] dout[0] dout[1] dout[2] dout[3] sram_rw_4bit
.ends sram_64x4_with_rw
** End of subcircuit definition.

** Cell name: adder_4bit_sign_extension
.subckt adder_4bit_sign_extension vdd gnd sign a[0] a[1] a[2] a[3] b[0] b[1] b[2] b[3] s[0] s[1] s[2] s[3] s[4] 
xi_ha_0 vdd gnd a[0] b[0] s[0] c[0] half_adder
xi_fa_1 vdd gnd a[1] b[1] c[0] s[1] c[1] full_adder
xi_fa_2 vdd gnd a[2] b[2] c[1] s[2] c[2] full_adder
xi_fa_3 vdd gnd a[3] b[3] c[2] s[3] c[3] full_adder
xi_fa_4 vdd gnd sign a[3] b[3] c[3] s[4] adder_sign_extension
.ends adder_4bit_sign_extension
** End of subcircuit definition.

** Cell name: adder_5bit_sign_extension
.subckt adder_5bit_sign_extension vdd gnd sign a[0] a[1] a[2] a[3] a[4] b[0] b[1] b[2] b[3] b[4] s[0] s[1] s[2] s[3] s[4] s[5] 
xi_ha_0 vdd gnd a[0] b[0] s[0] c[0] half_adder
xi_fa_1 vdd gnd a[1] b[1] c[0] s[1] c[1] full_adder
xi_fa_2 vdd gnd a[2] b[2] c[1] s[2] c[2] full_adder
xi_fa_3 vdd gnd a[3] b[3] c[2] s[3] c[3] full_adder
xi_fa_4 vdd gnd a[4] b[4] c[3] s[4] c[4] full_adder
xi_fa_5 vdd gnd sign a[4] b[4] c[4] s[5] adder_sign_extension
.ends adder_5bit_sign_extension
** End of subcircuit definition.

** Cell name: adder_6bit_sign_extension
.subckt adder_6bit_sign_extension vdd gnd sign a[0] a[1] a[2] a[3] a[4] a[5] b[0] b[1] b[2] b[3] b[4] b[5] s[0] s[1] s[2] s[3] s[4] s[5] s[6] 
xi_ha_0 vdd gnd a[0] b[0] s[0] c[0] half_adder
xi_fa_1 vdd gnd a[1] b[1] c[0] s[1] c[1] full_adder
xi_fa_2 vdd gnd a[2] b[2] c[1] s[2] c[2] full_adder
xi_fa_3 vdd gnd a[3] b[3] c[2] s[3] c[3] full_adder
xi_fa_4 vdd gnd a[4] b[4] c[3] s[4] c[4] full_adder
xi_fa_5 vdd gnd a[5] b[5] c[4] s[5] c[5] full_adder
xi_fa_6 vdd gnd sign a[5] b[5] c[5] s[6] adder_sign_extension
.ends adder_6bit_sign_extension
** End of subcircuit definition.

** Cell name: adder_7bit_sign_extension
.subckt adder_7bit_sign_extension vdd gnd sign a[0] a[1] a[2] a[3] a[4] a[5] a[6] b[0] b[1] b[2] b[3] b[4] b[5] b[6] s[0] s[1] s[2] s[3] s[4] s[5] s[6] s[7] 
xi_ha_0 vdd gnd a[0] b[0] s[0] c[0] half_adder
xi_fa_1 vdd gnd a[1] b[1] c[0] s[1] c[1] full_adder
xi_fa_2 vdd gnd a[2] b[2] c[1] s[2] c[2] full_adder
xi_fa_3 vdd gnd a[3] b[3] c[2] s[3] c[3] full_adder
xi_fa_4 vdd gnd a[4] b[4] c[3] s[4] c[4] full_adder
xi_fa_5 vdd gnd a[5] b[5] c[4] s[5] c[5] full_adder
xi_fa_6 vdd gnd a[6] b[6] c[5] s[6] c[6] full_adder
xi_fa_7 vdd gnd sign a[6] b[6] c[6] s[7] adder_sign_extension
.ends adder_7bit_sign_extension
** End of subcircuit definition.

** Cell name: adder_8bit_sign_extension
.subckt adder_8bit_sign_extension vdd gnd sign a[0] a[1] a[2] a[3] a[4] a[5] a[6] a[7] b[0] b[1] b[2] b[3] b[4] b[5] b[6] b[7] s[0] s[1] s[2] s[3] s[4] s[5] s[6] s[7] s[8] 
xi_ha_0 vdd gnd a[0] b[0] s[0] c[0] half_adder
xi_fa_1 vdd gnd a[1] b[1] c[0] s[1] c[1] full_adder
xi_fa_2 vdd gnd a[2] b[2] c[1] s[2] c[2] full_adder
xi_fa_3 vdd gnd a[3] b[3] c[2] s[3] c[3] full_adder
xi_fa_4 vdd gnd a[4] b[4] c[3] s[4] c[4] full_adder
xi_fa_5 vdd gnd a[5] b[5] c[4] s[5] c[5] full_adder
xi_fa_6 vdd gnd a[6] b[6] c[5] s[6] c[6] full_adder
xi_fa_7 vdd gnd a[7] b[7] c[6] s[7] c[7] full_adder
xi_fa_8 vdd gnd sign a[7] b[7] c[7] s[8] adder_sign_extension
.ends adder_8bit_sign_extension
** End of subcircuit definition.

** Cell name: adder_9bit_sign_extension
.subckt adder_9bit_sign_extension vdd gnd sign a[0] a[1] a[2] a[3] a[4] a[5] a[6] a[7] a[8] b[0] b[1] b[2] b[3] b[4] b[5] b[6] b[7] b[8] s[0] s[1] s[2] s[3] s[4] s[5] s[6] s[7] s[8] s[9] 
xi_ha_0 vdd gnd a[0] b[0] s[0] c[0] half_adder
xi_fa_1 vdd gnd a[1] b[1] c[0] s[1] c[1] full_adder
xi_fa_2 vdd gnd a[2] b[2] c[1] s[2] c[2] full_adder
xi_fa_3 vdd gnd a[3] b[3] c[2] s[3] c[3] full_adder
xi_fa_4 vdd gnd a[4] b[4] c[3] s[4] c[4] full_adder
xi_fa_5 vdd gnd a[5] b[5] c[4] s[5] c[5] full_adder
xi_fa_6 vdd gnd a[6] b[6] c[5] s[6] c[6] full_adder
xi_fa_7 vdd gnd a[7] b[7] c[6] s[7] c[7] full_adder
xi_fa_8 vdd gnd a[8] b[8] c[7] s[8] c[8] full_adder
xi_fa_9 vdd gnd sign a[8] b[8] c[8] s[9] adder_sign_extension
.ends adder_9bit_sign_extension
** End of subcircuit definition.

** Cell name: adder_tree_4bit_to_10bit
.subckt adder_tree_4bit_to_10bit vdd gnd sign_weight in_0[0] in_0[1] in_0[2] in_0[3] in_1[0] in_1[1] in_1[2] in_1[3] in_2[0] in_2[1] in_2[2] in_2[3] in_3[0] in_3[1] in_3[2] in_3[3] in_4[0] in_4[1] in_4[2] in_4[3] in_5[0] in_5[1] in_5[2] in_5[3] in_6[0] in_6[1] in_6[2] in_6[3] in_7[0] in_7[1] in_7[2] in_7[3] in_8[0] in_8[1] in_8[2] in_8[3] in_9[0] in_9[1] in_9[2] in_9[3] in_10[0] in_10[1] in_10[2] in_10[3] in_11[0] in_11[1] in_11[2] in_11[3] in_12[0] in_12[1] in_12[2] in_12[3] in_13[0] in_13[1] in_13[2] in_13[3] in_14[0] in_14[1] in_14[2] in_14[3] in_15[0] in_15[1] in_15[2] in_15[3] in_16[0] in_16[1] in_16[2] in_16[3] in_17[0] in_17[1] in_17[2] in_17[3] in_18[0] in_18[1] in_18[2] in_18[3] in_19[0] in_19[1] in_19[2] in_19[3] in_20[0] in_20[1] in_20[2] in_20[3] in_21[0] in_21[1] in_21[2] in_21[3] in_22[0] in_22[1] in_22[2] in_22[3] in_23[0] in_23[1] in_23[2] in_23[3] in_24[0] in_24[1] in_24[2] in_24[3] in_25[0] in_25[1] in_25[2] in_25[3] in_26[0] in_26[1] in_26[2] in_26[3] in_27[0] in_27[1] in_27[2] in_27[3] in_28[0] in_28[1] in_28[2] in_28[3] in_29[0] in_29[1] in_29[2] in_29[3] in_30[0] in_30[1] in_30[2] in_30[3] in_31[0] in_31[1] in_31[2] in_31[3] in_32[0] in_32[1] in_32[2] in_32[3] in_33[0] in_33[1] in_33[2] in_33[3] in_34[0] in_34[1] in_34[2] in_34[3] in_35[0] in_35[1] in_35[2] in_35[3] in_36[0] in_36[1] in_36[2] in_36[3] in_37[0] in_37[1] in_37[2] in_37[3] in_38[0] in_38[1] in_38[2] in_38[3] in_39[0] in_39[1] in_39[2] in_39[3] in_40[0] in_40[1] in_40[2] in_40[3] in_41[0] in_41[1] in_41[2] in_41[3] in_42[0] in_42[1] in_42[2] in_42[3] in_43[0] in_43[1] in_43[2] in_43[3] in_44[0] in_44[1] in_44[2] in_44[3] in_45[0] in_45[1] in_45[2] in_45[3] in_46[0] in_46[1] in_46[2] in_46[3] in_47[0] in_47[1] in_47[2] in_47[3] in_48[0] in_48[1] in_48[2] in_48[3] in_49[0] in_49[1] in_49[2] in_49[3] in_50[0] in_50[1] in_50[2] in_50[3] in_51[0] in_51[1] in_51[2] in_51[3] in_52[0] in_52[1] in_52[2] in_52[3] in_53[0] in_53[1] in_53[2] in_53[3] in_54[0] in_54[1] in_54[2] in_54[3] in_55[0] in_55[1] in_55[2] in_55[3] in_56[0] in_56[1] in_56[2] in_56[3] in_57[0] in_57[1] in_57[2] in_57[3] in_58[0] in_58[1] in_58[2] in_58[3] in_59[0] in_59[1] in_59[2] in_59[3] in_60[0] in_60[1] in_60[2] in_60[3] in_61[0] in_61[1] in_61[2] in_61[3] in_62[0] in_62[1] in_62[2] in_62[3] in_63[0] in_63[1] in_63[2] in_63[3] out[0] out[1] out[2] out[3] out[4] out[5] out[6] out[7] out[8] out[9] 
xi_adder_4bit_0 vdd gnd sign_weight in_0[0] in_0[1] in_0[2] in_0[3] in_1[0] in_1[1] in_1[2] in_1[3] sum_4bit_0[0] sum_4bit_0[1] sum_4bit_0[2] sum_4bit_0[3] sum_4bit_0[4] adder_4bit_sign_extension
xi_adder_4bit_1 vdd gnd sign_weight in_2[0] in_2[1] in_2[2] in_2[3] in_3[0] in_3[1] in_3[2] in_3[3] sum_4bit_1[0] sum_4bit_1[1] sum_4bit_1[2] sum_4bit_1[3] sum_4bit_1[4] adder_4bit_sign_extension
xi_adder_4bit_2 vdd gnd sign_weight in_4[0] in_4[1] in_4[2] in_4[3] in_5[0] in_5[1] in_5[2] in_5[3] sum_4bit_2[0] sum_4bit_2[1] sum_4bit_2[2] sum_4bit_2[3] sum_4bit_2[4] adder_4bit_sign_extension
xi_adder_4bit_3 vdd gnd sign_weight in_6[0] in_6[1] in_6[2] in_6[3] in_7[0] in_7[1] in_7[2] in_7[3] sum_4bit_3[0] sum_4bit_3[1] sum_4bit_3[2] sum_4bit_3[3] sum_4bit_3[4] adder_4bit_sign_extension
xi_adder_4bit_4 vdd gnd sign_weight in_8[0] in_8[1] in_8[2] in_8[3] in_9[0] in_9[1] in_9[2] in_9[3] sum_4bit_4[0] sum_4bit_4[1] sum_4bit_4[2] sum_4bit_4[3] sum_4bit_4[4] adder_4bit_sign_extension
xi_adder_4bit_5 vdd gnd sign_weight in_10[0] in_10[1] in_10[2] in_10[3] in_11[0] in_11[1] in_11[2] in_11[3] sum_4bit_5[0] sum_4bit_5[1] sum_4bit_5[2] sum_4bit_5[3] sum_4bit_5[4] adder_4bit_sign_extension
xi_adder_4bit_6 vdd gnd sign_weight in_12[0] in_12[1] in_12[2] in_12[3] in_13[0] in_13[1] in_13[2] in_13[3] sum_4bit_6[0] sum_4bit_6[1] sum_4bit_6[2] sum_4bit_6[3] sum_4bit_6[4] adder_4bit_sign_extension
xi_adder_4bit_7 vdd gnd sign_weight in_14[0] in_14[1] in_14[2] in_14[3] in_15[0] in_15[1] in_15[2] in_15[3] sum_4bit_7[0] sum_4bit_7[1] sum_4bit_7[2] sum_4bit_7[3] sum_4bit_7[4] adder_4bit_sign_extension
xi_adder_4bit_8 vdd gnd sign_weight in_16[0] in_16[1] in_16[2] in_16[3] in_17[0] in_17[1] in_17[2] in_17[3] sum_4bit_8[0] sum_4bit_8[1] sum_4bit_8[2] sum_4bit_8[3] sum_4bit_8[4] adder_4bit_sign_extension
xi_adder_4bit_9 vdd gnd sign_weight in_18[0] in_18[1] in_18[2] in_18[3] in_19[0] in_19[1] in_19[2] in_19[3] sum_4bit_9[0] sum_4bit_9[1] sum_4bit_9[2] sum_4bit_9[3] sum_4bit_9[4] adder_4bit_sign_extension
xi_adder_4bit_10 vdd gnd sign_weight in_20[0] in_20[1] in_20[2] in_20[3] in_21[0] in_21[1] in_21[2] in_21[3] sum_4bit_10[0] sum_4bit_10[1] sum_4bit_10[2] sum_4bit_10[3] sum_4bit_10[4] adder_4bit_sign_extension
xi_adder_4bit_11 vdd gnd sign_weight in_22[0] in_22[1] in_22[2] in_22[3] in_23[0] in_23[1] in_23[2] in_23[3] sum_4bit_11[0] sum_4bit_11[1] sum_4bit_11[2] sum_4bit_11[3] sum_4bit_11[4] adder_4bit_sign_extension
xi_adder_4bit_12 vdd gnd sign_weight in_24[0] in_24[1] in_24[2] in_24[3] in_25[0] in_25[1] in_25[2] in_25[3] sum_4bit_12[0] sum_4bit_12[1] sum_4bit_12[2] sum_4bit_12[3] sum_4bit_12[4] adder_4bit_sign_extension
xi_adder_4bit_13 vdd gnd sign_weight in_26[0] in_26[1] in_26[2] in_26[3] in_27[0] in_27[1] in_27[2] in_27[3] sum_4bit_13[0] sum_4bit_13[1] sum_4bit_13[2] sum_4bit_13[3] sum_4bit_13[4] adder_4bit_sign_extension
xi_adder_4bit_14 vdd gnd sign_weight in_28[0] in_28[1] in_28[2] in_28[3] in_29[0] in_29[1] in_29[2] in_29[3] sum_4bit_14[0] sum_4bit_14[1] sum_4bit_14[2] sum_4bit_14[3] sum_4bit_14[4] adder_4bit_sign_extension
xi_adder_4bit_15 vdd gnd sign_weight in_30[0] in_30[1] in_30[2] in_30[3] in_31[0] in_31[1] in_31[2] in_31[3] sum_4bit_15[0] sum_4bit_15[1] sum_4bit_15[2] sum_4bit_15[3] sum_4bit_15[4] adder_4bit_sign_extension
xi_adder_4bit_16 vdd gnd sign_weight in_32[0] in_32[1] in_32[2] in_32[3] in_33[0] in_33[1] in_33[2] in_33[3] sum_4bit_16[0] sum_4bit_16[1] sum_4bit_16[2] sum_4bit_16[3] sum_4bit_16[4] adder_4bit_sign_extension
xi_adder_4bit_17 vdd gnd sign_weight in_34[0] in_34[1] in_34[2] in_34[3] in_35[0] in_35[1] in_35[2] in_35[3] sum_4bit_17[0] sum_4bit_17[1] sum_4bit_17[2] sum_4bit_17[3] sum_4bit_17[4] adder_4bit_sign_extension
xi_adder_4bit_18 vdd gnd sign_weight in_36[0] in_36[1] in_36[2] in_36[3] in_37[0] in_37[1] in_37[2] in_37[3] sum_4bit_18[0] sum_4bit_18[1] sum_4bit_18[2] sum_4bit_18[3] sum_4bit_18[4] adder_4bit_sign_extension
xi_adder_4bit_19 vdd gnd sign_weight in_38[0] in_38[1] in_38[2] in_38[3] in_39[0] in_39[1] in_39[2] in_39[3] sum_4bit_19[0] sum_4bit_19[1] sum_4bit_19[2] sum_4bit_19[3] sum_4bit_19[4] adder_4bit_sign_extension
xi_adder_4bit_20 vdd gnd sign_weight in_40[0] in_40[1] in_40[2] in_40[3] in_41[0] in_41[1] in_41[2] in_41[3] sum_4bit_20[0] sum_4bit_20[1] sum_4bit_20[2] sum_4bit_20[3] sum_4bit_20[4] adder_4bit_sign_extension
xi_adder_4bit_21 vdd gnd sign_weight in_42[0] in_42[1] in_42[2] in_42[3] in_43[0] in_43[1] in_43[2] in_43[3] sum_4bit_21[0] sum_4bit_21[1] sum_4bit_21[2] sum_4bit_21[3] sum_4bit_21[4] adder_4bit_sign_extension
xi_adder_4bit_22 vdd gnd sign_weight in_44[0] in_44[1] in_44[2] in_44[3] in_45[0] in_45[1] in_45[2] in_45[3] sum_4bit_22[0] sum_4bit_22[1] sum_4bit_22[2] sum_4bit_22[3] sum_4bit_22[4] adder_4bit_sign_extension
xi_adder_4bit_23 vdd gnd sign_weight in_46[0] in_46[1] in_46[2] in_46[3] in_47[0] in_47[1] in_47[2] in_47[3] sum_4bit_23[0] sum_4bit_23[1] sum_4bit_23[2] sum_4bit_23[3] sum_4bit_23[4] adder_4bit_sign_extension
xi_adder_4bit_24 vdd gnd sign_weight in_48[0] in_48[1] in_48[2] in_48[3] in_49[0] in_49[1] in_49[2] in_49[3] sum_4bit_24[0] sum_4bit_24[1] sum_4bit_24[2] sum_4bit_24[3] sum_4bit_24[4] adder_4bit_sign_extension
xi_adder_4bit_25 vdd gnd sign_weight in_50[0] in_50[1] in_50[2] in_50[3] in_51[0] in_51[1] in_51[2] in_51[3] sum_4bit_25[0] sum_4bit_25[1] sum_4bit_25[2] sum_4bit_25[3] sum_4bit_25[4] adder_4bit_sign_extension
xi_adder_4bit_26 vdd gnd sign_weight in_52[0] in_52[1] in_52[2] in_52[3] in_53[0] in_53[1] in_53[2] in_53[3] sum_4bit_26[0] sum_4bit_26[1] sum_4bit_26[2] sum_4bit_26[3] sum_4bit_26[4] adder_4bit_sign_extension
xi_adder_4bit_27 vdd gnd sign_weight in_54[0] in_54[1] in_54[2] in_54[3] in_55[0] in_55[1] in_55[2] in_55[3] sum_4bit_27[0] sum_4bit_27[1] sum_4bit_27[2] sum_4bit_27[3] sum_4bit_27[4] adder_4bit_sign_extension
xi_adder_4bit_28 vdd gnd sign_weight in_56[0] in_56[1] in_56[2] in_56[3] in_57[0] in_57[1] in_57[2] in_57[3] sum_4bit_28[0] sum_4bit_28[1] sum_4bit_28[2] sum_4bit_28[3] sum_4bit_28[4] adder_4bit_sign_extension
xi_adder_4bit_29 vdd gnd sign_weight in_58[0] in_58[1] in_58[2] in_58[3] in_59[0] in_59[1] in_59[2] in_59[3] sum_4bit_29[0] sum_4bit_29[1] sum_4bit_29[2] sum_4bit_29[3] sum_4bit_29[4] adder_4bit_sign_extension
xi_adder_4bit_30 vdd gnd sign_weight in_60[0] in_60[1] in_60[2] in_60[3] in_61[0] in_61[1] in_61[2] in_61[3] sum_4bit_30[0] sum_4bit_30[1] sum_4bit_30[2] sum_4bit_30[3] sum_4bit_30[4] adder_4bit_sign_extension
xi_adder_4bit_31 vdd gnd sign_weight in_62[0] in_62[1] in_62[2] in_62[3] in_63[0] in_63[1] in_63[2] in_63[3] sum_4bit_31[0] sum_4bit_31[1] sum_4bit_31[2] sum_4bit_31[3] sum_4bit_31[4] adder_4bit_sign_extension
xi_adder_5bit_0 vdd gnd sign_weight sum_4bit_0[0] sum_4bit_0[1] sum_4bit_0[2] sum_4bit_0[3] sum_4bit_0[4] sum_4bit_1[0] sum_4bit_1[1] sum_4bit_1[2] sum_4bit_1[3] sum_4bit_1[4] sum_5bit_0[0] sum_5bit_0[1] sum_5bit_0[2] sum_5bit_0[3] sum_5bit_0[4] sum_5bit_0[5] adder_5bit_sign_extension
xi_adder_5bit_1 vdd gnd sign_weight sum_4bit_2[0] sum_4bit_2[1] sum_4bit_2[2] sum_4bit_2[3] sum_4bit_2[4] sum_4bit_3[0] sum_4bit_3[1] sum_4bit_3[2] sum_4bit_3[3] sum_4bit_3[4] sum_5bit_1[0] sum_5bit_1[1] sum_5bit_1[2] sum_5bit_1[3] sum_5bit_1[4] sum_5bit_1[5] adder_5bit_sign_extension
xi_adder_5bit_2 vdd gnd sign_weight sum_4bit_4[0] sum_4bit_4[1] sum_4bit_4[2] sum_4bit_4[3] sum_4bit_4[4] sum_4bit_5[0] sum_4bit_5[1] sum_4bit_5[2] sum_4bit_5[3] sum_4bit_5[4] sum_5bit_2[0] sum_5bit_2[1] sum_5bit_2[2] sum_5bit_2[3] sum_5bit_2[4] sum_5bit_2[5] adder_5bit_sign_extension
xi_adder_5bit_3 vdd gnd sign_weight sum_4bit_6[0] sum_4bit_6[1] sum_4bit_6[2] sum_4bit_6[3] sum_4bit_6[4] sum_4bit_7[0] sum_4bit_7[1] sum_4bit_7[2] sum_4bit_7[3] sum_4bit_7[4] sum_5bit_3[0] sum_5bit_3[1] sum_5bit_3[2] sum_5bit_3[3] sum_5bit_3[4] sum_5bit_3[5] adder_5bit_sign_extension
xi_adder_5bit_4 vdd gnd sign_weight sum_4bit_8[0] sum_4bit_8[1] sum_4bit_8[2] sum_4bit_8[3] sum_4bit_8[4] sum_4bit_9[0] sum_4bit_9[1] sum_4bit_9[2] sum_4bit_9[3] sum_4bit_9[4] sum_5bit_4[0] sum_5bit_4[1] sum_5bit_4[2] sum_5bit_4[3] sum_5bit_4[4] sum_5bit_4[5] adder_5bit_sign_extension
xi_adder_5bit_5 vdd gnd sign_weight sum_4bit_10[0] sum_4bit_10[1] sum_4bit_10[2] sum_4bit_10[3] sum_4bit_10[4] sum_4bit_11[0] sum_4bit_11[1] sum_4bit_11[2] sum_4bit_11[3] sum_4bit_11[4] sum_5bit_5[0] sum_5bit_5[1] sum_5bit_5[2] sum_5bit_5[3] sum_5bit_5[4] sum_5bit_5[5] adder_5bit_sign_extension
xi_adder_5bit_6 vdd gnd sign_weight sum_4bit_12[0] sum_4bit_12[1] sum_4bit_12[2] sum_4bit_12[3] sum_4bit_12[4] sum_4bit_13[0] sum_4bit_13[1] sum_4bit_13[2] sum_4bit_13[3] sum_4bit_13[4] sum_5bit_6[0] sum_5bit_6[1] sum_5bit_6[2] sum_5bit_6[3] sum_5bit_6[4] sum_5bit_6[5] adder_5bit_sign_extension
xi_adder_5bit_7 vdd gnd sign_weight sum_4bit_14[0] sum_4bit_14[1] sum_4bit_14[2] sum_4bit_14[3] sum_4bit_14[4] sum_4bit_15[0] sum_4bit_15[1] sum_4bit_15[2] sum_4bit_15[3] sum_4bit_15[4] sum_5bit_7[0] sum_5bit_7[1] sum_5bit_7[2] sum_5bit_7[3] sum_5bit_7[4] sum_5bit_7[5] adder_5bit_sign_extension
xi_adder_5bit_8 vdd gnd sign_weight sum_4bit_16[0] sum_4bit_16[1] sum_4bit_16[2] sum_4bit_16[3] sum_4bit_16[4] sum_4bit_17[0] sum_4bit_17[1] sum_4bit_17[2] sum_4bit_17[3] sum_4bit_17[4] sum_5bit_8[0] sum_5bit_8[1] sum_5bit_8[2] sum_5bit_8[3] sum_5bit_8[4] sum_5bit_8[5] adder_5bit_sign_extension
xi_adder_5bit_9 vdd gnd sign_weight sum_4bit_18[0] sum_4bit_18[1] sum_4bit_18[2] sum_4bit_18[3] sum_4bit_18[4] sum_4bit_19[0] sum_4bit_19[1] sum_4bit_19[2] sum_4bit_19[3] sum_4bit_19[4] sum_5bit_9[0] sum_5bit_9[1] sum_5bit_9[2] sum_5bit_9[3] sum_5bit_9[4] sum_5bit_9[5] adder_5bit_sign_extension
xi_adder_5bit_10 vdd gnd sign_weight sum_4bit_20[0] sum_4bit_20[1] sum_4bit_20[2] sum_4bit_20[3] sum_4bit_20[4] sum_4bit_21[0] sum_4bit_21[1] sum_4bit_21[2] sum_4bit_21[3] sum_4bit_21[4] sum_5bit_10[0] sum_5bit_10[1] sum_5bit_10[2] sum_5bit_10[3] sum_5bit_10[4] sum_5bit_10[5] adder_5bit_sign_extension
xi_adder_5bit_11 vdd gnd sign_weight sum_4bit_22[0] sum_4bit_22[1] sum_4bit_22[2] sum_4bit_22[3] sum_4bit_22[4] sum_4bit_23[0] sum_4bit_23[1] sum_4bit_23[2] sum_4bit_23[3] sum_4bit_23[4] sum_5bit_11[0] sum_5bit_11[1] sum_5bit_11[2] sum_5bit_11[3] sum_5bit_11[4] sum_5bit_11[5] adder_5bit_sign_extension
xi_adder_5bit_12 vdd gnd sign_weight sum_4bit_24[0] sum_4bit_24[1] sum_4bit_24[2] sum_4bit_24[3] sum_4bit_24[4] sum_4bit_25[0] sum_4bit_25[1] sum_4bit_25[2] sum_4bit_25[3] sum_4bit_25[4] sum_5bit_12[0] sum_5bit_12[1] sum_5bit_12[2] sum_5bit_12[3] sum_5bit_12[4] sum_5bit_12[5] adder_5bit_sign_extension
xi_adder_5bit_13 vdd gnd sign_weight sum_4bit_26[0] sum_4bit_26[1] sum_4bit_26[2] sum_4bit_26[3] sum_4bit_26[4] sum_4bit_27[0] sum_4bit_27[1] sum_4bit_27[2] sum_4bit_27[3] sum_4bit_27[4] sum_5bit_13[0] sum_5bit_13[1] sum_5bit_13[2] sum_5bit_13[3] sum_5bit_13[4] sum_5bit_13[5] adder_5bit_sign_extension
xi_adder_5bit_14 vdd gnd sign_weight sum_4bit_28[0] sum_4bit_28[1] sum_4bit_28[2] sum_4bit_28[3] sum_4bit_28[4] sum_4bit_29[0] sum_4bit_29[1] sum_4bit_29[2] sum_4bit_29[3] sum_4bit_29[4] sum_5bit_14[0] sum_5bit_14[1] sum_5bit_14[2] sum_5bit_14[3] sum_5bit_14[4] sum_5bit_14[5] adder_5bit_sign_extension
xi_adder_5bit_15 vdd gnd sign_weight sum_4bit_30[0] sum_4bit_30[1] sum_4bit_30[2] sum_4bit_30[3] sum_4bit_30[4] sum_4bit_31[0] sum_4bit_31[1] sum_4bit_31[2] sum_4bit_31[3] sum_4bit_31[4] sum_5bit_15[0] sum_5bit_15[1] sum_5bit_15[2] sum_5bit_15[3] sum_5bit_15[4] sum_5bit_15[5] adder_5bit_sign_extension
xi_adder_6bit_0 vdd gnd sign_weight sum_5bit_0[0] sum_5bit_0[1] sum_5bit_0[2] sum_5bit_0[3] sum_5bit_0[4] sum_5bit_0[5] sum_5bit_1[0] sum_5bit_1[1] sum_5bit_1[2] sum_5bit_1[3] sum_5bit_1[4] sum_5bit_1[5] sum_6bit_0[0] sum_6bit_0[1] sum_6bit_0[2] sum_6bit_0[3] sum_6bit_0[4] sum_6bit_0[5] sum_6bit_0[6] adder_6bit_sign_extension
xi_adder_6bit_1 vdd gnd sign_weight sum_5bit_2[0] sum_5bit_2[1] sum_5bit_2[2] sum_5bit_2[3] sum_5bit_2[4] sum_5bit_2[5] sum_5bit_3[0] sum_5bit_3[1] sum_5bit_3[2] sum_5bit_3[3] sum_5bit_3[4] sum_5bit_3[5] sum_6bit_1[0] sum_6bit_1[1] sum_6bit_1[2] sum_6bit_1[3] sum_6bit_1[4] sum_6bit_1[5] sum_6bit_1[6] adder_6bit_sign_extension
xi_adder_6bit_2 vdd gnd sign_weight sum_5bit_4[0] sum_5bit_4[1] sum_5bit_4[2] sum_5bit_4[3] sum_5bit_4[4] sum_5bit_4[5] sum_5bit_5[0] sum_5bit_5[1] sum_5bit_5[2] sum_5bit_5[3] sum_5bit_5[4] sum_5bit_5[5] sum_6bit_2[0] sum_6bit_2[1] sum_6bit_2[2] sum_6bit_2[3] sum_6bit_2[4] sum_6bit_2[5] sum_6bit_2[6] adder_6bit_sign_extension
xi_adder_6bit_3 vdd gnd sign_weight sum_5bit_6[0] sum_5bit_6[1] sum_5bit_6[2] sum_5bit_6[3] sum_5bit_6[4] sum_5bit_6[5] sum_5bit_7[0] sum_5bit_7[1] sum_5bit_7[2] sum_5bit_7[3] sum_5bit_7[4] sum_5bit_7[5] sum_6bit_3[0] sum_6bit_3[1] sum_6bit_3[2] sum_6bit_3[3] sum_6bit_3[4] sum_6bit_3[5] sum_6bit_3[6] adder_6bit_sign_extension
xi_adder_6bit_4 vdd gnd sign_weight sum_5bit_8[0] sum_5bit_8[1] sum_5bit_8[2] sum_5bit_8[3] sum_5bit_8[4] sum_5bit_8[5] sum_5bit_9[0] sum_5bit_9[1] sum_5bit_9[2] sum_5bit_9[3] sum_5bit_9[4] sum_5bit_9[5] sum_6bit_4[0] sum_6bit_4[1] sum_6bit_4[2] sum_6bit_4[3] sum_6bit_4[4] sum_6bit_4[5] sum_6bit_4[6] adder_6bit_sign_extension
xi_adder_6bit_5 vdd gnd sign_weight sum_5bit_10[0] sum_5bit_10[1] sum_5bit_10[2] sum_5bit_10[3] sum_5bit_10[4] sum_5bit_10[5] sum_5bit_11[0] sum_5bit_11[1] sum_5bit_11[2] sum_5bit_11[3] sum_5bit_11[4] sum_5bit_11[5] sum_6bit_5[0] sum_6bit_5[1] sum_6bit_5[2] sum_6bit_5[3] sum_6bit_5[4] sum_6bit_5[5] sum_6bit_5[6] adder_6bit_sign_extension
xi_adder_6bit_6 vdd gnd sign_weight sum_5bit_12[0] sum_5bit_12[1] sum_5bit_12[2] sum_5bit_12[3] sum_5bit_12[4] sum_5bit_12[5] sum_5bit_13[0] sum_5bit_13[1] sum_5bit_13[2] sum_5bit_13[3] sum_5bit_13[4] sum_5bit_13[5] sum_6bit_6[0] sum_6bit_6[1] sum_6bit_6[2] sum_6bit_6[3] sum_6bit_6[4] sum_6bit_6[5] sum_6bit_6[6] adder_6bit_sign_extension
xi_adder_6bit_7 vdd gnd sign_weight sum_5bit_14[0] sum_5bit_14[1] sum_5bit_14[2] sum_5bit_14[3] sum_5bit_14[4] sum_5bit_14[5] sum_5bit_15[0] sum_5bit_15[1] sum_5bit_15[2] sum_5bit_15[3] sum_5bit_15[4] sum_5bit_15[5] sum_6bit_7[0] sum_6bit_7[1] sum_6bit_7[2] sum_6bit_7[3] sum_6bit_7[4] sum_6bit_7[5] sum_6bit_7[6] adder_6bit_sign_extension
xi_adder_7bit_0 vdd gnd sign_weight sum_6bit_0[0] sum_6bit_0[1] sum_6bit_0[2] sum_6bit_0[3] sum_6bit_0[4] sum_6bit_0[5] sum_6bit_0[6] sum_6bit_1[0] sum_6bit_1[1] sum_6bit_1[2] sum_6bit_1[3] sum_6bit_1[4] sum_6bit_1[5] sum_6bit_1[6] sum_7bit_0[0] sum_7bit_0[1] sum_7bit_0[2] sum_7bit_0[3] sum_7bit_0[4] sum_7bit_0[5] sum_7bit_0[6] sum_7bit_0[7] adder_7bit_sign_extension
xi_adder_7bit_1 vdd gnd sign_weight sum_6bit_2[0] sum_6bit_2[1] sum_6bit_2[2] sum_6bit_2[3] sum_6bit_2[4] sum_6bit_2[5] sum_6bit_2[6] sum_6bit_3[0] sum_6bit_3[1] sum_6bit_3[2] sum_6bit_3[3] sum_6bit_3[4] sum_6bit_3[5] sum_6bit_3[6] sum_7bit_1[0] sum_7bit_1[1] sum_7bit_1[2] sum_7bit_1[3] sum_7bit_1[4] sum_7bit_1[5] sum_7bit_1[6] sum_7bit_1[7] adder_7bit_sign_extension
xi_adder_7bit_2 vdd gnd sign_weight sum_6bit_4[0] sum_6bit_4[1] sum_6bit_4[2] sum_6bit_4[3] sum_6bit_4[4] sum_6bit_4[5] sum_6bit_4[6] sum_6bit_5[0] sum_6bit_5[1] sum_6bit_5[2] sum_6bit_5[3] sum_6bit_5[4] sum_6bit_5[5] sum_6bit_5[6] sum_7bit_2[0] sum_7bit_2[1] sum_7bit_2[2] sum_7bit_2[3] sum_7bit_2[4] sum_7bit_2[5] sum_7bit_2[6] sum_7bit_2[7] adder_7bit_sign_extension
xi_adder_7bit_3 vdd gnd sign_weight sum_6bit_6[0] sum_6bit_6[1] sum_6bit_6[2] sum_6bit_6[3] sum_6bit_6[4] sum_6bit_6[5] sum_6bit_6[6] sum_6bit_7[0] sum_6bit_7[1] sum_6bit_7[2] sum_6bit_7[3] sum_6bit_7[4] sum_6bit_7[5] sum_6bit_7[6] sum_7bit_3[0] sum_7bit_3[1] sum_7bit_3[2] sum_7bit_3[3] sum_7bit_3[4] sum_7bit_3[5] sum_7bit_3[6] sum_7bit_3[7] adder_7bit_sign_extension
xi_adder_8bit_0 vdd gnd sign_weight sum_7bit_0[0] sum_7bit_0[1] sum_7bit_0[2] sum_7bit_0[3] sum_7bit_0[4] sum_7bit_0[5] sum_7bit_0[6] sum_7bit_0[7] sum_7bit_1[0] sum_7bit_1[1] sum_7bit_1[2] sum_7bit_1[3] sum_7bit_1[4] sum_7bit_1[5] sum_7bit_1[6] sum_7bit_1[7] sum_8bit_0[0] sum_8bit_0[1] sum_8bit_0[2] sum_8bit_0[3] sum_8bit_0[4] sum_8bit_0[5] sum_8bit_0[6] sum_8bit_0[7] sum_8bit_0[8] adder_8bit_sign_extension
xi_adder_8bit_1 vdd gnd sign_weight sum_7bit_2[0] sum_7bit_2[1] sum_7bit_2[2] sum_7bit_2[3] sum_7bit_2[4] sum_7bit_2[5] sum_7bit_2[6] sum_7bit_2[7] sum_7bit_3[0] sum_7bit_3[1] sum_7bit_3[2] sum_7bit_3[3] sum_7bit_3[4] sum_7bit_3[5] sum_7bit_3[6] sum_7bit_3[7] sum_8bit_1[0] sum_8bit_1[1] sum_8bit_1[2] sum_8bit_1[3] sum_8bit_1[4] sum_8bit_1[5] sum_8bit_1[6] sum_8bit_1[7] sum_8bit_1[8] adder_8bit_sign_extension
xi_adder_9bit vdd gnd sign_weight sum_8bit_0[0] sum_8bit_0[1] sum_8bit_0[2] sum_8bit_0[3] sum_8bit_0[4] sum_8bit_0[5] sum_8bit_0[6] sum_8bit_0[7] sum_8bit_0[8] sum_8bit_1[0] sum_8bit_1[1] sum_8bit_1[2] sum_8bit_1[3] sum_8bit_1[4] sum_8bit_1[5] sum_8bit_1[6] sum_8bit_1[7] sum_8bit_1[8] out[0] out[1] out[2] out[3] out[4] out[5] out[6] out[7] out[8] out[9] adder_9bit_sign_extension
.ends adder_tree_4bit_to_10bit
** End of subcircuit definition.

** Cell name: adder_14bit_with_cin_for_acc
.subckt adder_14bit_with_cin_for_acc vdd gnd c_in a_0_to_9[0] a_0_to_9[1] a_0_to_9[2] a_0_to_9[3] a_0_to_9[4] a_0_to_9[5] a_0_to_9[6] a_0_to_9[7] a_0_to_9[8] a_0_to_9[9] a_10 a_11 a_12 a_13 b_0 b_1_to_13[0] b_1_to_13[1] b_1_to_13[2] b_1_to_13[3] b_1_to_13[4] b_1_to_13[5] b_1_to_13[6] b_1_to_13[7] b_1_to_13[8] b_1_to_13[9] b_1_to_13[10] b_1_to_13[11] b_1_to_13[12] s[0] s[1] s[2] s[3] s[4] s[5] s[6] s[7] s[8] s[9] s[10] s[11] s[12] s[13] 
xi_fa_0 vdd gnd a_0_to_9[0] b_0 c_in s[0] c[0] full_adder
xi_fa_1 vdd gnd a_0_to_9[1] b_1_to_13[0] c[0] s[1] c[1] full_adder
xi_fa_2 vdd gnd a_0_to_9[2] b_1_to_13[1] c[1] s[2] c[2] full_adder
xi_fa_3 vdd gnd a_0_to_9[3] b_1_to_13[2] c[2] s[3] c[3] full_adder
xi_fa_4 vdd gnd a_0_to_9[4] b_1_to_13[3] c[3] s[4] c[4] full_adder
xi_fa_5 vdd gnd a_0_to_9[5] b_1_to_13[4] c[4] s[5] c[5] full_adder
xi_fa_6 vdd gnd a_0_to_9[6] b_1_to_13[5] c[5] s[6] c[6] full_adder
xi_fa_7 vdd gnd a_0_to_9[7] b_1_to_13[6] c[6] s[7] c[7] full_adder
xi_fa_8 vdd gnd a_0_to_9[8] b_1_to_13[7] c[7] s[8] c[8] full_adder
xi_fa_9 vdd gnd a_0_to_9[9] b_1_to_13[8] c[8] s[9] c[9] full_adder
xi_fa_10 vdd gnd a_10 b_1_to_13[9] c[9] s[10] c[10] full_adder
xi_fa_11 vdd gnd a_11 b_1_to_13[10] c[10] s[11] c[11] full_adder
xi_fa_12 vdd gnd a_12 b_1_to_13[11] c[11] s[12] c[12] full_adder
xi_fa_13 vdd gnd a_13 b_1_to_13[12] c[12] s[13] c[13] full_adder
.ends adder_14bit_with_cin_for_acc
** End of subcircuit definition.

** Cell name: dff_10bit
.subckt dff_10bit vdd gnd clk rst_b in[0] in[1] in[2] in[3] in[4] in[5] in[6] in[7] in[8] in[9] out[0] out[1] out[2] out[3] out[4] out[5] out[6] out[7] out[8] out[9] 
xi_dff_0 vdd gnd clk rst_b in_0 out_0 dff
xi_dff_1 vdd gnd clk rst_b in_1 out_1 dff
xi_dff_2 vdd gnd clk rst_b in_2 out_2 dff
xi_dff_3 vdd gnd clk rst_b in_3 out_3 dff
xi_dff_4 vdd gnd clk rst_b in_4 out_4 dff
xi_dff_5 vdd gnd clk rst_b in_5 out_5 dff
xi_dff_6 vdd gnd clk rst_b in_6 out_6 dff
xi_dff_7 vdd gnd clk rst_b in_7 out_7 dff
xi_dff_8 vdd gnd clk rst_b in_8 out_8 dff
xi_dff_9 vdd gnd clk rst_b in_9 out_9 dff
.ends dff_10bit
** End of subcircuit definition.

** Cell name: dff_13bit
.subckt dff_13bit vdd gnd clk rst_b in[0] in[1] in[2] in[3] in[4] in[5] in[6] in[7] in[8] in[9] in[10] in[11] in[12] out[0] out[1] out[2] out[3] out[4] out[5] out[6] out[7] out[8] out[9] out[10] out[11] out[12] 
xi_dff_0 vdd gnd clk rst_b in_0 out_0 dff
xi_dff_1 vdd gnd clk rst_b in_1 out_1 dff
xi_dff_2 vdd gnd clk rst_b in_2 out_2 dff
xi_dff_3 vdd gnd clk rst_b in_3 out_3 dff
xi_dff_4 vdd gnd clk rst_b in_4 out_4 dff
xi_dff_5 vdd gnd clk rst_b in_5 out_5 dff
xi_dff_6 vdd gnd clk rst_b in_6 out_6 dff
xi_dff_7 vdd gnd clk rst_b in_7 out_7 dff
xi_dff_8 vdd gnd clk rst_b in_8 out_8 dff
xi_dff_9 vdd gnd clk rst_b in_9 out_9 dff
xi_dff_10 vdd gnd clk rst_b in_10 out_10 dff
xi_dff_11 vdd gnd clk rst_b in_11 out_11 dff
xi_dff_12 vdd gnd clk rst_b in_12 out_12 dff
.ends dff_13bit
** End of subcircuit definition.

** Cell name: dff_14bit
.subckt dff_14bit vdd gnd clk rst_b in[0] in[1] in[2] in[3] in[4] in[5] in[6] in[7] in[8] in[9] in[10] in[11] in[12] in[13] out[0] out[1] out[2] out[3] out[4] out[5] out[6] out[7] out[8] out[9] out[10] out[11] out[12] out[13] 
xi_dff_0 vdd gnd clk rst_b in_0 out_0 dff
xi_dff_1 vdd gnd clk rst_b in_1 out_1 dff
xi_dff_2 vdd gnd clk rst_b in_2 out_2 dff
xi_dff_3 vdd gnd clk rst_b in_3 out_3 dff
xi_dff_4 vdd gnd clk rst_b in_4 out_4 dff
xi_dff_5 vdd gnd clk rst_b in_5 out_5 dff
xi_dff_6 vdd gnd clk rst_b in_6 out_6 dff
xi_dff_7 vdd gnd clk rst_b in_7 out_7 dff
xi_dff_8 vdd gnd clk rst_b in_8 out_8 dff
xi_dff_9 vdd gnd clk rst_b in_9 out_9 dff
xi_dff_10 vdd gnd clk rst_b in_10 out_10 dff
xi_dff_11 vdd gnd clk rst_b in_11 out_11 dff
xi_dff_12 vdd gnd clk rst_b in_12 out_12 dff
xi_dff_13 vdd gnd clk rst_b in_13 out_13 dff
.ends dff_14bit
** End of subcircuit definition.

** Cell name: inverse_mux_10bit
.subckt inverse_mux_10bit sign vdd gnd in[0] in[1] in[2] in[3] in[4] in[5] in[6] in[7] in[8] in[9] out[0] out[1] out[2] out[3] out[4] out[5] out[6] out[7] out[8] out[9] 
xi_inv_sign vdd gnd sign sign_b inverter
xi_inv_in_0 vdd gnd in[0] in_b[0] inverter
xi_inv_in_1 vdd gnd in[1] in_b[1] inverter
xi_inv_in_2 vdd gnd in[2] in_b[2] inverter
xi_inv_in_3 vdd gnd in[3] in_b[3] inverter
xi_inv_in_4 vdd gnd in[4] in_b[4] inverter
xi_inv_in_5 vdd gnd in[5] in_b[5] inverter
xi_inv_in_6 vdd gnd in[6] in_b[6] inverter
xi_inv_in_7 vdd gnd in[7] in_b[7] inverter
xi_inv_in_8 vdd gnd in[8] in_b[8] inverter
xi_inv_in_9 vdd gnd in[9] in_b[9] inverter
xi_in_0_0 vdd gnd in[0] sign_b in_0[0] nand2
xi_in_1_0 vdd gnd in_b[0] sign in_1[0] nand2
xi_in_0_1 vdd gnd in[1] sign_b in_0[1] nand2
xi_in_1_1 vdd gnd in_b[1] sign in_1[1] nand2
xi_in_0_2 vdd gnd in[2] sign_b in_0[2] nand2
xi_in_1_2 vdd gnd in_b[2] sign in_1[2] nand2
xi_in_0_3 vdd gnd in[3] sign_b in_0[3] nand2
xi_in_1_3 vdd gnd in_b[3] sign in_1[3] nand2
xi_in_0_4 vdd gnd in[4] sign_b in_0[4] nand2
xi_in_1_4 vdd gnd in_b[4] sign in_1[4] nand2
xi_in_0_5 vdd gnd in[5] sign_b in_0[5] nand2
xi_in_1_5 vdd gnd in_b[5] sign in_1[5] nand2
xi_in_0_6 vdd gnd in[6] sign_b in_0[6] nand2
xi_in_1_6 vdd gnd in_b[6] sign in_1[6] nand2
xi_in_0_7 vdd gnd in[7] sign_b in_0[7] nand2
xi_in_1_7 vdd gnd in_b[7] sign in_1[7] nand2
xi_in_0_8 vdd gnd in[8] sign_b in_0[8] nand2
xi_in_1_8 vdd gnd in_b[8] sign in_1[8] nand2
xi_in_0_9 vdd gnd in[9] sign_b in_0[9] nand2
xi_in_1_9 vdd gnd in_b[9] sign in_1[9] nand2
xi_out_0 vdd gnd in_0[0] in_1[0] out[0] nand2
xi_out_1 vdd gnd in_0[1] in_1[1] out[1] nand2
xi_out_2 vdd gnd in_0[2] in_1[2] out[2] nand2
xi_out_3 vdd gnd in_0[3] in_1[3] out[3] nand2
xi_out_4 vdd gnd in_0[4] in_1[4] out[4] nand2
xi_out_5 vdd gnd in_0[5] in_1[5] out[5] nand2
xi_out_6 vdd gnd in_0[6] in_1[6] out[6] nand2
xi_out_7 vdd gnd in_0[7] in_1[7] out[7] nand2
xi_out_8 vdd gnd in_0[8] in_1[8] out[8] nand2
xi_out_9 vdd gnd in_0[9] in_1[9] out[9] nand2
.ends inverse_mux_10bit
** End of subcircuit definition.

** Cell name: accumulator_10bit_to_14bit
.subckt accumulator_10bit_to_14bit vdd gnd clk_psum clk_shift clk_out rst_b_psum rst_b_shift rst_b_out sign_weight sign_in in_msb in[0] in[1] in[2] in[3] in[4] in[5] in[6] in[7] in[8] in[9] out[0] out[1] out[2] out[3] out[4] out[5] out[6] out[7] out[8] out[9] out[10] out[11] out[12] out[13] 
xi_dff_psum vdd gnd clk_psum rst_b_psum in[0] in[1] in[2] in[3] in[4] in[5] in[6] in[7] in[8] in[9] psum[0] psum[1] psum[2] psum[3] psum[4] psum[5] psum[6] psum[7] psum[8] psum[9] dff_10bit
xi_nand_acc vdd gnd sign_in in_msb sign_in_msb_b nand2
xi_inv_acc vdd gnd sign_in_msb_b sign_in_msb inverter
xi_inverse_mux vdd gnd sign_in_msb psum[0] psum[1] psum[2] psum[3] psum[4] psum[5] psum[6] psum[7] psum[8] psum[9] complement[0] complement[1] complement[2] complement[3] complement[4] complement[5] complement[6] complement[7] complement[8] complement[9] inverse_mux_10bit
xi_mux vdd gnd sign_weight sign_in_msb complement[9] extension mux_2_1
xi_adder vdd gnd sign_in_msb complement[0] complement[1] complement[2] complement[3] complement[4] complement[5] complement[6] complement[7] complement[8] complement[9] extension extension extension extension gnd shift[0] shift[1] shift[2] shift[3] shift[4] shift[5] shift[6] shift[7] shift[8] shift[9] shift[10] shift[11] shift[12] sum[0] sum[1] sum[2] sum[3] sum[4] sum[5] sum[6] sum[7] sum[8] sum[9] sum[10] sum[11] sum[12] sum[13] adder_14bit_with_cin_for_acc
xi_dff_shift vdd gnd clk_shift rst_b_shift sum[0] sum[1] sum[2] sum[3] sum[4] sum[5] sum[6] sum[7] sum[8] sum[9] sum[10] sum[11] sum[12] shift[0] shift[1] shift[2] shift[3] shift[4] shift[5] shift[6] shift[7] shift[8] shift[9] shift[10] shift[11] shift[12] dff_13bit
xi_dff_out vdd gnd clk_out rst_b_out sum[0] sum[1] sum[2] sum[3] sum[4] sum[5] sum[6] sum[7] sum[8] sum[9] sum[10] sum[11] sum[12] sum[13] out[0] out[1] out[2] out[3] out[4] out[5] out[6] out[7] out[8] out[9] out[10] out[11] out[12] out[13] dff_14bit
.ends accumulator_10bit_to_14bit
** End of subcircuit definition.

** Cell name: dcim_column_64x4x4
.subckt dcim_column_64x4x4 vdd gnd clk_psum clk_shift clk_out rst_b_psum rst_b_shift rst_b_out sign_weight sign_in in_msb pe ysw ysr spe se wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] in_b[0] in_b[1] in_b[2] in_b[3] in_b[4] in_b[5] in_b[6] in_b[7] in_b[8] in_b[9] in_b[10] in_b[11] in_b[12] in_b[13] in_b[14] in_b[15] in_b[16] in_b[17] in_b[18] in_b[19] in_b[20] in_b[21] in_b[22] in_b[23] in_b[24] in_b[25] in_b[26] in_b[27] in_b[28] in_b[29] in_b[30] in_b[31] in_b[32] in_b[33] in_b[34] in_b[35] in_b[36] in_b[37] in_b[38] in_b[39] in_b[40] in_b[41] in_b[42] in_b[43] in_b[44] in_b[45] in_b[46] in_b[47] in_b[48] in_b[49] in_b[50] in_b[51] in_b[52] in_b[53] in_b[54] in_b[55] in_b[56] in_b[57] in_b[58] in_b[59] in_b[60] in_b[61] in_b[62] in_b[63] din[0] din[1] din[2] din[3] dout[0] dout[1] dout[2] dout[3] column_psum[0] column_psum[1] column_psum[2] column_psum[3] column_psum[4] column_psum[5] column_psum[6] column_psum[7] column_psum[8] column_psum[9] column_psum[10] column_psum[11] column_psum[12] column_psum[13] 
xi_sram_with_rw vdd gnd pe ysw ysr spe se wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] in_b[0] in_b[1] in_b[2] in_b[3] in_b[4] in_b[5] in_b[6] in_b[7] in_b[8] in_b[9] in_b[10] in_b[11] in_b[12] in_b[13] in_b[14] in_b[15] in_b[16] in_b[17] in_b[18] in_b[19] in_b[20] in_b[21] in_b[22] in_b[23] in_b[24] in_b[25] in_b[26] in_b[27] in_b[28] in_b[29] in_b[30] in_b[31] in_b[32] in_b[33] in_b[34] in_b[35] in_b[36] in_b[37] in_b[38] in_b[39] in_b[40] in_b[41] in_b[42] in_b[43] in_b[44] in_b[45] in_b[46] in_b[47] in_b[48] in_b[49] in_b[50] in_b[51] in_b[52] in_b[53] in_b[54] in_b[55] in_b[56] in_b[57] in_b[58] in_b[59] in_b[60] in_b[61] in_b[62] in_b[63] din[0] din[1] din[2] din[3] dout[0] dout[1] dout[2] dout[3] bitcell_out_0[0] bitcell_out_0[1] bitcell_out_0[2] bitcell_out_0[3] bitcell_out_1[0] bitcell_out_1[1] bitcell_out_1[2] bitcell_out_1[3] bitcell_out_2[0] bitcell_out_2[1] bitcell_out_2[2] bitcell_out_2[3] bitcell_out_3[0] bitcell_out_3[1] bitcell_out_3[2] bitcell_out_3[3] bitcell_out_4[0] bitcell_out_4[1] bitcell_out_4[2] bitcell_out_4[3] bitcell_out_5[0] bitcell_out_5[1] bitcell_out_5[2] bitcell_out_5[3] bitcell_out_6[0] bitcell_out_6[1] bitcell_out_6[2] bitcell_out_6[3] bitcell_out_7[0] bitcell_out_7[1] bitcell_out_7[2] bitcell_out_7[3] bitcell_out_8[0] bitcell_out_8[1] bitcell_out_8[2] bitcell_out_8[3] bitcell_out_9[0] bitcell_out_9[1] bitcell_out_9[2] bitcell_out_9[3] bitcell_out_10[0] bitcell_out_10[1] bitcell_out_10[2] bitcell_out_10[3] bitcell_out_11[0] bitcell_out_11[1] bitcell_out_11[2] bitcell_out_11[3] bitcell_out_12[0] bitcell_out_12[1] bitcell_out_12[2] bitcell_out_12[3] bitcell_out_13[0] bitcell_out_13[1] bitcell_out_13[2] bitcell_out_13[3] bitcell_out_14[0] bitcell_out_14[1] bitcell_out_14[2] bitcell_out_14[3] bitcell_out_15[0] bitcell_out_15[1] bitcell_out_15[2] bitcell_out_15[3] bitcell_out_16[0] bitcell_out_16[1] bitcell_out_16[2] bitcell_out_16[3] bitcell_out_17[0] bitcell_out_17[1] bitcell_out_17[2] bitcell_out_17[3] bitcell_out_18[0] bitcell_out_18[1] bitcell_out_18[2] bitcell_out_18[3] bitcell_out_19[0] bitcell_out_19[1] bitcell_out_19[2] bitcell_out_19[3] bitcell_out_20[0] bitcell_out_20[1] bitcell_out_20[2] bitcell_out_20[3] bitcell_out_21[0] bitcell_out_21[1] bitcell_out_21[2] bitcell_out_21[3] bitcell_out_22[0] bitcell_out_22[1] bitcell_out_22[2] bitcell_out_22[3] bitcell_out_23[0] bitcell_out_23[1] bitcell_out_23[2] bitcell_out_23[3] bitcell_out_24[0] bitcell_out_24[1] bitcell_out_24[2] bitcell_out_24[3] bitcell_out_25[0] bitcell_out_25[1] bitcell_out_25[2] bitcell_out_25[3] bitcell_out_26[0] bitcell_out_26[1] bitcell_out_26[2] bitcell_out_26[3] bitcell_out_27[0] bitcell_out_27[1] bitcell_out_27[2] bitcell_out_27[3] bitcell_out_28[0] bitcell_out_28[1] bitcell_out_28[2] bitcell_out_28[3] bitcell_out_29[0] bitcell_out_29[1] bitcell_out_29[2] bitcell_out_29[3] bitcell_out_30[0] bitcell_out_30[1] bitcell_out_30[2] bitcell_out_30[3] bitcell_out_31[0] bitcell_out_31[1] bitcell_out_31[2] bitcell_out_31[3] bitcell_out_32[0] bitcell_out_32[1] bitcell_out_32[2] bitcell_out_32[3] bitcell_out_33[0] bitcell_out_33[1] bitcell_out_33[2] bitcell_out_33[3] bitcell_out_34[0] bitcell_out_34[1] bitcell_out_34[2] bitcell_out_34[3] bitcell_out_35[0] bitcell_out_35[1] bitcell_out_35[2] bitcell_out_35[3] bitcell_out_36[0] bitcell_out_36[1] bitcell_out_36[2] bitcell_out_36[3] bitcell_out_37[0] bitcell_out_37[1] bitcell_out_37[2] bitcell_out_37[3] bitcell_out_38[0] bitcell_out_38[1] bitcell_out_38[2] bitcell_out_38[3] bitcell_out_39[0] bitcell_out_39[1] bitcell_out_39[2] bitcell_out_39[3] bitcell_out_40[0] bitcell_out_40[1] bitcell_out_40[2] bitcell_out_40[3] bitcell_out_41[0] bitcell_out_41[1] bitcell_out_41[2] bitcell_out_41[3] bitcell_out_42[0] bitcell_out_42[1] bitcell_out_42[2] bitcell_out_42[3] bitcell_out_43[0] bitcell_out_43[1] bitcell_out_43[2] bitcell_out_43[3] bitcell_out_44[0] bitcell_out_44[1] bitcell_out_44[2] bitcell_out_44[3] bitcell_out_45[0] bitcell_out_45[1] bitcell_out_45[2] bitcell_out_45[3] bitcell_out_46[0] bitcell_out_46[1] bitcell_out_46[2] bitcell_out_46[3] bitcell_out_47[0] bitcell_out_47[1] bitcell_out_47[2] bitcell_out_47[3] bitcell_out_48[0] bitcell_out_48[1] bitcell_out_48[2] bitcell_out_48[3] bitcell_out_49[0] bitcell_out_49[1] bitcell_out_49[2] bitcell_out_49[3] bitcell_out_50[0] bitcell_out_50[1] bitcell_out_50[2] bitcell_out_50[3] bitcell_out_51[0] bitcell_out_51[1] bitcell_out_51[2] bitcell_out_51[3] bitcell_out_52[0] bitcell_out_52[1] bitcell_out_52[2] bitcell_out_52[3] bitcell_out_53[0] bitcell_out_53[1] bitcell_out_53[2] bitcell_out_53[3] bitcell_out_54[0] bitcell_out_54[1] bitcell_out_54[2] bitcell_out_54[3] bitcell_out_55[0] bitcell_out_55[1] bitcell_out_55[2] bitcell_out_55[3] bitcell_out_56[0] bitcell_out_56[1] bitcell_out_56[2] bitcell_out_56[3] bitcell_out_57[0] bitcell_out_57[1] bitcell_out_57[2] bitcell_out_57[3] bitcell_out_58[0] bitcell_out_58[1] bitcell_out_58[2] bitcell_out_58[3] bitcell_out_59[0] bitcell_out_59[1] bitcell_out_59[2] bitcell_out_59[3] bitcell_out_60[0] bitcell_out_60[1] bitcell_out_60[2] bitcell_out_60[3] bitcell_out_61[0] bitcell_out_61[1] bitcell_out_61[2] bitcell_out_61[3] bitcell_out_62[0] bitcell_out_62[1] bitcell_out_62[2] bitcell_out_62[3] bitcell_out_63[0] bitcell_out_63[1] bitcell_out_63[2] bitcell_out_63[3] sram_64x4_with_rw
xi_adder_tree vdd gnd sign_weight bitcell_out_0[0] bitcell_out_0[1] bitcell_out_0[2] bitcell_out_0[3] bitcell_out_1[0] bitcell_out_1[1] bitcell_out_1[2] bitcell_out_1[3] bitcell_out_2[0] bitcell_out_2[1] bitcell_out_2[2] bitcell_out_2[3] bitcell_out_3[0] bitcell_out_3[1] bitcell_out_3[2] bitcell_out_3[3] bitcell_out_4[0] bitcell_out_4[1] bitcell_out_4[2] bitcell_out_4[3] bitcell_out_5[0] bitcell_out_5[1] bitcell_out_5[2] bitcell_out_5[3] bitcell_out_6[0] bitcell_out_6[1] bitcell_out_6[2] bitcell_out_6[3] bitcell_out_7[0] bitcell_out_7[1] bitcell_out_7[2] bitcell_out_7[3] bitcell_out_8[0] bitcell_out_8[1] bitcell_out_8[2] bitcell_out_8[3] bitcell_out_9[0] bitcell_out_9[1] bitcell_out_9[2] bitcell_out_9[3] bitcell_out_10[0] bitcell_out_10[1] bitcell_out_10[2] bitcell_out_10[3] bitcell_out_11[0] bitcell_out_11[1] bitcell_out_11[2] bitcell_out_11[3] bitcell_out_12[0] bitcell_out_12[1] bitcell_out_12[2] bitcell_out_12[3] bitcell_out_13[0] bitcell_out_13[1] bitcell_out_13[2] bitcell_out_13[3] bitcell_out_14[0] bitcell_out_14[1] bitcell_out_14[2] bitcell_out_14[3] bitcell_out_15[0] bitcell_out_15[1] bitcell_out_15[2] bitcell_out_15[3] bitcell_out_16[0] bitcell_out_16[1] bitcell_out_16[2] bitcell_out_16[3] bitcell_out_17[0] bitcell_out_17[1] bitcell_out_17[2] bitcell_out_17[3] bitcell_out_18[0] bitcell_out_18[1] bitcell_out_18[2] bitcell_out_18[3] bitcell_out_19[0] bitcell_out_19[1] bitcell_out_19[2] bitcell_out_19[3] bitcell_out_20[0] bitcell_out_20[1] bitcell_out_20[2] bitcell_out_20[3] bitcell_out_21[0] bitcell_out_21[1] bitcell_out_21[2] bitcell_out_21[3] bitcell_out_22[0] bitcell_out_22[1] bitcell_out_22[2] bitcell_out_22[3] bitcell_out_23[0] bitcell_out_23[1] bitcell_out_23[2] bitcell_out_23[3] bitcell_out_24[0] bitcell_out_24[1] bitcell_out_24[2] bitcell_out_24[3] bitcell_out_25[0] bitcell_out_25[1] bitcell_out_25[2] bitcell_out_25[3] bitcell_out_26[0] bitcell_out_26[1] bitcell_out_26[2] bitcell_out_26[3] bitcell_out_27[0] bitcell_out_27[1] bitcell_out_27[2] bitcell_out_27[3] bitcell_out_28[0] bitcell_out_28[1] bitcell_out_28[2] bitcell_out_28[3] bitcell_out_29[0] bitcell_out_29[1] bitcell_out_29[2] bitcell_out_29[3] bitcell_out_30[0] bitcell_out_30[1] bitcell_out_30[2] bitcell_out_30[3] bitcell_out_31[0] bitcell_out_31[1] bitcell_out_31[2] bitcell_out_31[3] bitcell_out_32[0] bitcell_out_32[1] bitcell_out_32[2] bitcell_out_32[3] bitcell_out_33[0] bitcell_out_33[1] bitcell_out_33[2] bitcell_out_33[3] bitcell_out_34[0] bitcell_out_34[1] bitcell_out_34[2] bitcell_out_34[3] bitcell_out_35[0] bitcell_out_35[1] bitcell_out_35[2] bitcell_out_35[3] bitcell_out_36[0] bitcell_out_36[1] bitcell_out_36[2] bitcell_out_36[3] bitcell_out_37[0] bitcell_out_37[1] bitcell_out_37[2] bitcell_out_37[3] bitcell_out_38[0] bitcell_out_38[1] bitcell_out_38[2] bitcell_out_38[3] bitcell_out_39[0] bitcell_out_39[1] bitcell_out_39[2] bitcell_out_39[3] bitcell_out_40[0] bitcell_out_40[1] bitcell_out_40[2] bitcell_out_40[3] bitcell_out_41[0] bitcell_out_41[1] bitcell_out_41[2] bitcell_out_41[3] bitcell_out_42[0] bitcell_out_42[1] bitcell_out_42[2] bitcell_out_42[3] bitcell_out_43[0] bitcell_out_43[1] bitcell_out_43[2] bitcell_out_43[3] bitcell_out_44[0] bitcell_out_44[1] bitcell_out_44[2] bitcell_out_44[3] bitcell_out_45[0] bitcell_out_45[1] bitcell_out_45[2] bitcell_out_45[3] bitcell_out_46[0] bitcell_out_46[1] bitcell_out_46[2] bitcell_out_46[3] bitcell_out_47[0] bitcell_out_47[1] bitcell_out_47[2] bitcell_out_47[3] bitcell_out_48[0] bitcell_out_48[1] bitcell_out_48[2] bitcell_out_48[3] bitcell_out_49[0] bitcell_out_49[1] bitcell_out_49[2] bitcell_out_49[3] bitcell_out_50[0] bitcell_out_50[1] bitcell_out_50[2] bitcell_out_50[3] bitcell_out_51[0] bitcell_out_51[1] bitcell_out_51[2] bitcell_out_51[3] bitcell_out_52[0] bitcell_out_52[1] bitcell_out_52[2] bitcell_out_52[3] bitcell_out_53[0] bitcell_out_53[1] bitcell_out_53[2] bitcell_out_53[3] bitcell_out_54[0] bitcell_out_54[1] bitcell_out_54[2] bitcell_out_54[3] bitcell_out_55[0] bitcell_out_55[1] bitcell_out_55[2] bitcell_out_55[3] bitcell_out_56[0] bitcell_out_56[1] bitcell_out_56[2] bitcell_out_56[3] bitcell_out_57[0] bitcell_out_57[1] bitcell_out_57[2] bitcell_out_57[3] bitcell_out_58[0] bitcell_out_58[1] bitcell_out_58[2] bitcell_out_58[3] bitcell_out_59[0] bitcell_out_59[1] bitcell_out_59[2] bitcell_out_59[3] bitcell_out_60[0] bitcell_out_60[1] bitcell_out_60[2] bitcell_out_60[3] bitcell_out_61[0] bitcell_out_61[1] bitcell_out_61[2] bitcell_out_61[3] bitcell_out_62[0] bitcell_out_62[1] bitcell_out_62[2] bitcell_out_62[3] bitcell_out_63[0] bitcell_out_63[1] bitcell_out_63[2] bitcell_out_63[3] psum[0] psum[1] psum[2] psum[3] psum[4] psum[5] psum[6] psum[7] psum[8] psum[9] adder_tree_4bit_to_10bit
xi_accumulator vdd gnd clk_psum clk_shift clk_out rst_b_psum rst_b_shift rst_b_out sign_weight sign_in, in_msb psum[0] psum[1] psum[2] psum[3] psum[4] psum[5] psum[6] psum[7] psum[8] psum[9] column_psum[0] column_psum[1] column_psum[2] column_psum[3] column_psum[4] column_psum[5] column_psum[6] column_psum[7] column_psum[8] column_psum[9] column_psum[10] column_psum[11] column_psum[12] column_psum[13] accumulator_10bit_to_14bit
.ends dcim_column_64x4x4
** End of subcircuit definition.

