
module driver_64x64(\in<0> , \in<1> , \in<2> , \in<3> , \in<4> , \in<5> , \in<6> , \in<7> , \in<8> , \in<9> , \in<10> , \in<11> , \in<12> , \in<13> , \in<14> , \in<15> , \in<16> , \in<17> , \in<18> , \in<19> , \in<20> , \in<21> , \in<22> , \in<23> , \in<24> , \in<25> , \in<26> , \in<27> , \in<28> , \in<29> , \in<30> , \in<31> , \in<32> , \in<33> , \in<34> , \in<35> , \in<36> , \in<37> , \in<38> , \in<39> , \in<40> , \in<41> , \in<42> , \in<43> , \in<44> , \in<45> , \in<46> , \in<47> , \in<48> , \in<49> , \in<50> , \in<51> , \in<52> , \in<53> , \in<54> , \in<55> , \in<56> , \in<57> , \in<58> , \in<59> , \in<60> , \in<61> , \in<62> , \in<63> , \out<0> , \out<1> , \out<2> , \out<3> , \out<4> , \out<5> , \out<6> , \out<7> , \out<8> , \out<9> , \out<10> , \out<11> , \out<12> , \out<13> , \out<14> , \out<15> , \out<16> , \out<17> , \out<18> , \out<19> , \out<20> , \out<21> , \out<22> , \out<23> , \out<24> , \out<25> , \out<26> , \out<27> , \out<28> , \out<29> , \out<30> , \out<31> , \out<32> , \out<33> , \out<34> , \out<35> , \out<36> , \out<37> , \out<38> , \out<39> , \out<40> , \out<41> , \out<42> , \out<43> , \out<44> , \out<45> , \out<46> , \out<47> , \out<48> , \out<49> , \out<50> , \out<51> , \out<52> , \out<53> , \out<54> , \out<55> , \out<56> , \out<57> , \out<58> , \out<59> , \out<60> , \out<61> , \out<62> , \out<63> );
  input \in<0> ;
  input \in<10> ;
  input \in<11> ;
  input \in<12> ;
  input \in<13> ;
  input \in<14> ;
  input \in<15> ;
  input \in<16> ;
  input \in<17> ;
  input \in<18> ;
  input \in<19> ;
  input \in<1> ;
  input \in<20> ;
  input \in<21> ;
  input \in<22> ;
  input \in<23> ;
  input \in<24> ;
  input \in<25> ;
  input \in<26> ;
  input \in<27> ;
  input \in<28> ;
  input \in<29> ;
  input \in<2> ;
  input \in<30> ;
  input \in<31> ;
  input \in<32> ;
  input \in<33> ;
  input \in<34> ;
  input \in<35> ;
  input \in<36> ;
  input \in<37> ;
  input \in<38> ;
  input \in<39> ;
  input \in<3> ;
  input \in<40> ;
  input \in<41> ;
  input \in<42> ;
  input \in<43> ;
  input \in<44> ;
  input \in<45> ;
  input \in<46> ;
  input \in<47> ;
  input \in<48> ;
  input \in<49> ;
  input \in<4> ;
  input \in<50> ;
  input \in<51> ;
  input \in<52> ;
  input \in<53> ;
  input \in<54> ;
  input \in<55> ;
  input \in<56> ;
  input \in<57> ;
  input \in<58> ;
  input \in<59> ;
  input \in<5> ;
  input \in<60> ;
  input \in<61> ;
  input \in<62> ;
  input \in<63> ;
  input \in<6> ;
  input \in<7> ;
  input \in<8> ;
  input \in<9> ;
  wire \inv4_stage1_0.in ;
  wire \inv4_stage1_0.out ;
  wire \inv4_stage1_1.in ;
  wire \inv4_stage1_1.out ;
  wire \inv4_stage1_10.in ;
  wire \inv4_stage1_10.out ;
  wire \inv4_stage1_11.in ;
  wire \inv4_stage1_11.out ;
  wire \inv4_stage1_12.in ;
  wire \inv4_stage1_12.out ;
  wire \inv4_stage1_13.in ;
  wire \inv4_stage1_13.out ;
  wire \inv4_stage1_14.in ;
  wire \inv4_stage1_14.out ;
  wire \inv4_stage1_15.in ;
  wire \inv4_stage1_15.out ;
  wire \inv4_stage1_16.in ;
  wire \inv4_stage1_16.out ;
  wire \inv4_stage1_17.in ;
  wire \inv4_stage1_17.out ;
  wire \inv4_stage1_18.in ;
  wire \inv4_stage1_18.out ;
  wire \inv4_stage1_19.in ;
  wire \inv4_stage1_19.out ;
  wire \inv4_stage1_2.in ;
  wire \inv4_stage1_2.out ;
  wire \inv4_stage1_20.in ;
  wire \inv4_stage1_20.out ;
  wire \inv4_stage1_21.in ;
  wire \inv4_stage1_21.out ;
  wire \inv4_stage1_22.in ;
  wire \inv4_stage1_22.out ;
  wire \inv4_stage1_23.in ;
  wire \inv4_stage1_23.out ;
  wire \inv4_stage1_24.in ;
  wire \inv4_stage1_24.out ;
  wire \inv4_stage1_25.in ;
  wire \inv4_stage1_25.out ;
  wire \inv4_stage1_26.in ;
  wire \inv4_stage1_26.out ;
  wire \inv4_stage1_27.in ;
  wire \inv4_stage1_27.out ;
  wire \inv4_stage1_28.in ;
  wire \inv4_stage1_28.out ;
  wire \inv4_stage1_29.in ;
  wire \inv4_stage1_29.out ;
  wire \inv4_stage1_3.in ;
  wire \inv4_stage1_3.out ;
  wire \inv4_stage1_30.in ;
  wire \inv4_stage1_30.out ;
  wire \inv4_stage1_31.in ;
  wire \inv4_stage1_31.out ;
  wire \inv4_stage1_32.in ;
  wire \inv4_stage1_32.out ;
  wire \inv4_stage1_33.in ;
  wire \inv4_stage1_33.out ;
  wire \inv4_stage1_34.in ;
  wire \inv4_stage1_34.out ;
  wire \inv4_stage1_35.in ;
  wire \inv4_stage1_35.out ;
  wire \inv4_stage1_36.in ;
  wire \inv4_stage1_36.out ;
  wire \inv4_stage1_37.in ;
  wire \inv4_stage1_37.out ;
  wire \inv4_stage1_38.in ;
  wire \inv4_stage1_38.out ;
  wire \inv4_stage1_39.in ;
  wire \inv4_stage1_39.out ;
  wire \inv4_stage1_4.in ;
  wire \inv4_stage1_4.out ;
  wire \inv4_stage1_40.in ;
  wire \inv4_stage1_40.out ;
  wire \inv4_stage1_41.in ;
  wire \inv4_stage1_41.out ;
  wire \inv4_stage1_42.in ;
  wire \inv4_stage1_42.out ;
  wire \inv4_stage1_43.in ;
  wire \inv4_stage1_43.out ;
  wire \inv4_stage1_44.in ;
  wire \inv4_stage1_44.out ;
  wire \inv4_stage1_45.in ;
  wire \inv4_stage1_45.out ;
  wire \inv4_stage1_46.in ;
  wire \inv4_stage1_46.out ;
  wire \inv4_stage1_47.in ;
  wire \inv4_stage1_47.out ;
  wire \inv4_stage1_48.in ;
  wire \inv4_stage1_48.out ;
  wire \inv4_stage1_49.in ;
  wire \inv4_stage1_49.out ;
  wire \inv4_stage1_5.in ;
  wire \inv4_stage1_5.out ;
  wire \inv4_stage1_50.in ;
  wire \inv4_stage1_50.out ;
  wire \inv4_stage1_51.in ;
  wire \inv4_stage1_51.out ;
  wire \inv4_stage1_52.in ;
  wire \inv4_stage1_52.out ;
  wire \inv4_stage1_53.in ;
  wire \inv4_stage1_53.out ;
  wire \inv4_stage1_54.in ;
  wire \inv4_stage1_54.out ;
  wire \inv4_stage1_55.in ;
  wire \inv4_stage1_55.out ;
  wire \inv4_stage1_56.in ;
  wire \inv4_stage1_56.out ;
  wire \inv4_stage1_57.in ;
  wire \inv4_stage1_57.out ;
  wire \inv4_stage1_58.in ;
  wire \inv4_stage1_58.out ;
  wire \inv4_stage1_59.in ;
  wire \inv4_stage1_59.out ;
  wire \inv4_stage1_6.in ;
  wire \inv4_stage1_6.out ;
  wire \inv4_stage1_60.in ;
  wire \inv4_stage1_60.out ;
  wire \inv4_stage1_61.in ;
  wire \inv4_stage1_61.out ;
  wire \inv4_stage1_62.in ;
  wire \inv4_stage1_62.out ;
  wire \inv4_stage1_63.in ;
  wire \inv4_stage1_63.out ;
  wire \inv4_stage1_7.in ;
  wire \inv4_stage1_7.out ;
  wire \inv4_stage1_8.in ;
  wire \inv4_stage1_8.out ;
  wire \inv4_stage1_9.in ;
  wire \inv4_stage1_9.out ;
  output \out<0> ;
  output \out<10> ;
  output \out<11> ;
  output \out<12> ;
  output \out<13> ;
  output \out<14> ;
  output \out<15> ;
  output \out<16> ;
  output \out<17> ;
  output \out<18> ;
  output \out<19> ;
  output \out<1> ;
  output \out<20> ;
  output \out<21> ;
  output \out<22> ;
  output \out<23> ;
  output \out<24> ;
  output \out<25> ;
  output \out<26> ;
  output \out<27> ;
  output \out<28> ;
  output \out<29> ;
  output \out<2> ;
  output \out<30> ;
  output \out<31> ;
  output \out<32> ;
  output \out<33> ;
  output \out<34> ;
  output \out<35> ;
  output \out<36> ;
  output \out<37> ;
  output \out<38> ;
  output \out<39> ;
  output \out<3> ;
  output \out<40> ;
  output \out<41> ;
  output \out<42> ;
  output \out<43> ;
  output \out<44> ;
  output \out<45> ;
  output \out<46> ;
  output \out<47> ;
  output \out<48> ;
  output \out<49> ;
  output \out<4> ;
  output \out<50> ;
  output \out<51> ;
  output \out<52> ;
  output \out<53> ;
  output \out<54> ;
  output \out<55> ;
  output \out<56> ;
  output \out<57> ;
  output \out<58> ;
  output \out<59> ;
  output \out<5> ;
  output \out<60> ;
  output \out<61> ;
  output \out<62> ;
  output \out<63> ;
  output \out<6> ;
  output \out<7> ;
  output \out<8> ;
  output \out<9> ;
  wire \out_b<0> ;
  wire \out_b<10> ;
  wire \out_b<11> ;
  wire \out_b<12> ;
  wire \out_b<13> ;
  wire \out_b<14> ;
  wire \out_b<15> ;
  wire \out_b<16> ;
  wire \out_b<17> ;
  wire \out_b<18> ;
  wire \out_b<19> ;
  wire \out_b<1> ;
  wire \out_b<20> ;
  wire \out_b<21> ;
  wire \out_b<22> ;
  wire \out_b<23> ;
  wire \out_b<24> ;
  wire \out_b<25> ;
  wire \out_b<26> ;
  wire \out_b<27> ;
  wire \out_b<28> ;
  wire \out_b<29> ;
  wire \out_b<2> ;
  wire \out_b<30> ;
  wire \out_b<31> ;
  wire \out_b<32> ;
  wire \out_b<33> ;
  wire \out_b<34> ;
  wire \out_b<35> ;
  wire \out_b<36> ;
  wire \out_b<37> ;
  wire \out_b<38> ;
  wire \out_b<39> ;
  wire \out_b<3> ;
  wire \out_b<40> ;
  wire \out_b<41> ;
  wire \out_b<42> ;
  wire \out_b<43> ;
  wire \out_b<44> ;
  wire \out_b<45> ;
  wire \out_b<46> ;
  wire \out_b<47> ;
  wire \out_b<48> ;
  wire \out_b<49> ;
  wire \out_b<4> ;
  wire \out_b<50> ;
  wire \out_b<51> ;
  wire \out_b<52> ;
  wire \out_b<53> ;
  wire \out_b<54> ;
  wire \out_b<55> ;
  wire \out_b<56> ;
  wire \out_b<57> ;
  wire \out_b<58> ;
  wire \out_b<59> ;
  wire \out_b<5> ;
  wire \out_b<60> ;
  wire \out_b<61> ;
  wire \out_b<62> ;
  wire \out_b<63> ;
  wire \out_b<6> ;
  wire \out_b<7> ;
  wire \out_b<8> ;
  wire \out_b<9> ;
  inverter \inv4_stage1_0.inv_0  (    .in(\inv4_stage1_0.in ),    .out(\inv4_stage1_0.out )
  );
  inverter \inv4_stage1_0.inv_1  (    .in(\inv4_stage1_0.in ),    .out(\inv4_stage1_0.out )
  );
  inverter \inv4_stage1_0.inv_2  (    .in(\inv4_stage1_0.in ),    .out(\inv4_stage1_0.out )
  );
  inverter \inv4_stage1_0.inv_3  (    .in(\inv4_stage1_0.in ),    .out(\inv4_stage1_0.out )
  );
  inverter \inv4_stage1_1.inv_0  (    .in(\inv4_stage1_1.in ),    .out(\inv4_stage1_1.out )
  );
  inverter \inv4_stage1_1.inv_1  (    .in(\inv4_stage1_1.in ),    .out(\inv4_stage1_1.out )
  );
  inverter \inv4_stage1_1.inv_2  (    .in(\inv4_stage1_1.in ),    .out(\inv4_stage1_1.out )
  );
  inverter \inv4_stage1_1.inv_3  (    .in(\inv4_stage1_1.in ),    .out(\inv4_stage1_1.out )
  );
  inverter \inv4_stage1_10.inv_0  (    .in(\inv4_stage1_10.in ),    .out(\inv4_stage1_10.out )
  );
  inverter \inv4_stage1_10.inv_1  (    .in(\inv4_stage1_10.in ),    .out(\inv4_stage1_10.out )
  );
  inverter \inv4_stage1_10.inv_2  (    .in(\inv4_stage1_10.in ),    .out(\inv4_stage1_10.out )
  );
  inverter \inv4_stage1_10.inv_3  (    .in(\inv4_stage1_10.in ),    .out(\inv4_stage1_10.out )
  );
  inverter \inv4_stage1_11.inv_0  (    .in(\inv4_stage1_11.in ),    .out(\inv4_stage1_11.out )
  );
  inverter \inv4_stage1_11.inv_1  (    .in(\inv4_stage1_11.in ),    .out(\inv4_stage1_11.out )
  );
  inverter \inv4_stage1_11.inv_2  (    .in(\inv4_stage1_11.in ),    .out(\inv4_stage1_11.out )
  );
  inverter \inv4_stage1_11.inv_3  (    .in(\inv4_stage1_11.in ),    .out(\inv4_stage1_11.out )
  );
  inverter \inv4_stage1_12.inv_0  (    .in(\inv4_stage1_12.in ),    .out(\inv4_stage1_12.out )
  );
  inverter \inv4_stage1_12.inv_1  (    .in(\inv4_stage1_12.in ),    .out(\inv4_stage1_12.out )
  );
  inverter \inv4_stage1_12.inv_2  (    .in(\inv4_stage1_12.in ),    .out(\inv4_stage1_12.out )
  );
  inverter \inv4_stage1_12.inv_3  (    .in(\inv4_stage1_12.in ),    .out(\inv4_stage1_12.out )
  );
  inverter \inv4_stage1_13.inv_0  (    .in(\inv4_stage1_13.in ),    .out(\inv4_stage1_13.out )
  );
  inverter \inv4_stage1_13.inv_1  (    .in(\inv4_stage1_13.in ),    .out(\inv4_stage1_13.out )
  );
  inverter \inv4_stage1_13.inv_2  (    .in(\inv4_stage1_13.in ),    .out(\inv4_stage1_13.out )
  );
  inverter \inv4_stage1_13.inv_3  (    .in(\inv4_stage1_13.in ),    .out(\inv4_stage1_13.out )
  );
  inverter \inv4_stage1_14.inv_0  (    .in(\inv4_stage1_14.in ),    .out(\inv4_stage1_14.out )
  );
  inverter \inv4_stage1_14.inv_1  (    .in(\inv4_stage1_14.in ),    .out(\inv4_stage1_14.out )
  );
  inverter \inv4_stage1_14.inv_2  (    .in(\inv4_stage1_14.in ),    .out(\inv4_stage1_14.out )
  );
  inverter \inv4_stage1_14.inv_3  (    .in(\inv4_stage1_14.in ),    .out(\inv4_stage1_14.out )
  );
  inverter \inv4_stage1_15.inv_0  (    .in(\inv4_stage1_15.in ),    .out(\inv4_stage1_15.out )
  );
  inverter \inv4_stage1_15.inv_1  (    .in(\inv4_stage1_15.in ),    .out(\inv4_stage1_15.out )
  );
  inverter \inv4_stage1_15.inv_2  (    .in(\inv4_stage1_15.in ),    .out(\inv4_stage1_15.out )
  );
  inverter \inv4_stage1_15.inv_3  (    .in(\inv4_stage1_15.in ),    .out(\inv4_stage1_15.out )
  );
  inverter \inv4_stage1_16.inv_0  (    .in(\inv4_stage1_16.in ),    .out(\inv4_stage1_16.out )
  );
  inverter \inv4_stage1_16.inv_1  (    .in(\inv4_stage1_16.in ),    .out(\inv4_stage1_16.out )
  );
  inverter \inv4_stage1_16.inv_2  (    .in(\inv4_stage1_16.in ),    .out(\inv4_stage1_16.out )
  );
  inverter \inv4_stage1_16.inv_3  (    .in(\inv4_stage1_16.in ),    .out(\inv4_stage1_16.out )
  );
  inverter \inv4_stage1_17.inv_0  (    .in(\inv4_stage1_17.in ),    .out(\inv4_stage1_17.out )
  );
  inverter \inv4_stage1_17.inv_1  (    .in(\inv4_stage1_17.in ),    .out(\inv4_stage1_17.out )
  );
  inverter \inv4_stage1_17.inv_2  (    .in(\inv4_stage1_17.in ),    .out(\inv4_stage1_17.out )
  );
  inverter \inv4_stage1_17.inv_3  (    .in(\inv4_stage1_17.in ),    .out(\inv4_stage1_17.out )
  );
  inverter \inv4_stage1_18.inv_0  (    .in(\inv4_stage1_18.in ),    .out(\inv4_stage1_18.out )
  );
  inverter \inv4_stage1_18.inv_1  (    .in(\inv4_stage1_18.in ),    .out(\inv4_stage1_18.out )
  );
  inverter \inv4_stage1_18.inv_2  (    .in(\inv4_stage1_18.in ),    .out(\inv4_stage1_18.out )
  );
  inverter \inv4_stage1_18.inv_3  (    .in(\inv4_stage1_18.in ),    .out(\inv4_stage1_18.out )
  );
  inverter \inv4_stage1_19.inv_0  (    .in(\inv4_stage1_19.in ),    .out(\inv4_stage1_19.out )
  );
  inverter \inv4_stage1_19.inv_1  (    .in(\inv4_stage1_19.in ),    .out(\inv4_stage1_19.out )
  );
  inverter \inv4_stage1_19.inv_2  (    .in(\inv4_stage1_19.in ),    .out(\inv4_stage1_19.out )
  );
  inverter \inv4_stage1_19.inv_3  (    .in(\inv4_stage1_19.in ),    .out(\inv4_stage1_19.out )
  );
  inverter \inv4_stage1_2.inv_0  (    .in(\inv4_stage1_2.in ),    .out(\inv4_stage1_2.out )
  );
  inverter \inv4_stage1_2.inv_1  (    .in(\inv4_stage1_2.in ),    .out(\inv4_stage1_2.out )
  );
  inverter \inv4_stage1_2.inv_2  (    .in(\inv4_stage1_2.in ),    .out(\inv4_stage1_2.out )
  );
  inverter \inv4_stage1_2.inv_3  (    .in(\inv4_stage1_2.in ),    .out(\inv4_stage1_2.out )
  );
  inverter \inv4_stage1_20.inv_0  (    .in(\inv4_stage1_20.in ),    .out(\inv4_stage1_20.out )
  );
  inverter \inv4_stage1_20.inv_1  (    .in(\inv4_stage1_20.in ),    .out(\inv4_stage1_20.out )
  );
  inverter \inv4_stage1_20.inv_2  (    .in(\inv4_stage1_20.in ),    .out(\inv4_stage1_20.out )
  );
  inverter \inv4_stage1_20.inv_3  (    .in(\inv4_stage1_20.in ),    .out(\inv4_stage1_20.out )
  );
  inverter \inv4_stage1_21.inv_0  (    .in(\inv4_stage1_21.in ),    .out(\inv4_stage1_21.out )
  );
  inverter \inv4_stage1_21.inv_1  (    .in(\inv4_stage1_21.in ),    .out(\inv4_stage1_21.out )
  );
  inverter \inv4_stage1_21.inv_2  (    .in(\inv4_stage1_21.in ),    .out(\inv4_stage1_21.out )
  );
  inverter \inv4_stage1_21.inv_3  (    .in(\inv4_stage1_21.in ),    .out(\inv4_stage1_21.out )
  );
  inverter \inv4_stage1_22.inv_0  (    .in(\inv4_stage1_22.in ),    .out(\inv4_stage1_22.out )
  );
  inverter \inv4_stage1_22.inv_1  (    .in(\inv4_stage1_22.in ),    .out(\inv4_stage1_22.out )
  );
  inverter \inv4_stage1_22.inv_2  (    .in(\inv4_stage1_22.in ),    .out(\inv4_stage1_22.out )
  );
  inverter \inv4_stage1_22.inv_3  (    .in(\inv4_stage1_22.in ),    .out(\inv4_stage1_22.out )
  );
  inverter \inv4_stage1_23.inv_0  (    .in(\inv4_stage1_23.in ),    .out(\inv4_stage1_23.out )
  );
  inverter \inv4_stage1_23.inv_1  (    .in(\inv4_stage1_23.in ),    .out(\inv4_stage1_23.out )
  );
  inverter \inv4_stage1_23.inv_2  (    .in(\inv4_stage1_23.in ),    .out(\inv4_stage1_23.out )
  );
  inverter \inv4_stage1_23.inv_3  (    .in(\inv4_stage1_23.in ),    .out(\inv4_stage1_23.out )
  );
  inverter \inv4_stage1_24.inv_0  (    .in(\inv4_stage1_24.in ),    .out(\inv4_stage1_24.out )
  );
  inverter \inv4_stage1_24.inv_1  (    .in(\inv4_stage1_24.in ),    .out(\inv4_stage1_24.out )
  );
  inverter \inv4_stage1_24.inv_2  (    .in(\inv4_stage1_24.in ),    .out(\inv4_stage1_24.out )
  );
  inverter \inv4_stage1_24.inv_3  (    .in(\inv4_stage1_24.in ),    .out(\inv4_stage1_24.out )
  );
  inverter \inv4_stage1_25.inv_0  (    .in(\inv4_stage1_25.in ),    .out(\inv4_stage1_25.out )
  );
  inverter \inv4_stage1_25.inv_1  (    .in(\inv4_stage1_25.in ),    .out(\inv4_stage1_25.out )
  );
  inverter \inv4_stage1_25.inv_2  (    .in(\inv4_stage1_25.in ),    .out(\inv4_stage1_25.out )
  );
  inverter \inv4_stage1_25.inv_3  (    .in(\inv4_stage1_25.in ),    .out(\inv4_stage1_25.out )
  );
  inverter \inv4_stage1_26.inv_0  (    .in(\inv4_stage1_26.in ),    .out(\inv4_stage1_26.out )
  );
  inverter \inv4_stage1_26.inv_1  (    .in(\inv4_stage1_26.in ),    .out(\inv4_stage1_26.out )
  );
  inverter \inv4_stage1_26.inv_2  (    .in(\inv4_stage1_26.in ),    .out(\inv4_stage1_26.out )
  );
  inverter \inv4_stage1_26.inv_3  (    .in(\inv4_stage1_26.in ),    .out(\inv4_stage1_26.out )
  );
  inverter \inv4_stage1_27.inv_0  (    .in(\inv4_stage1_27.in ),    .out(\inv4_stage1_27.out )
  );
  inverter \inv4_stage1_27.inv_1  (    .in(\inv4_stage1_27.in ),    .out(\inv4_stage1_27.out )
  );
  inverter \inv4_stage1_27.inv_2  (    .in(\inv4_stage1_27.in ),    .out(\inv4_stage1_27.out )
  );
  inverter \inv4_stage1_27.inv_3  (    .in(\inv4_stage1_27.in ),    .out(\inv4_stage1_27.out )
  );
  inverter \inv4_stage1_28.inv_0  (    .in(\inv4_stage1_28.in ),    .out(\inv4_stage1_28.out )
  );
  inverter \inv4_stage1_28.inv_1  (    .in(\inv4_stage1_28.in ),    .out(\inv4_stage1_28.out )
  );
  inverter \inv4_stage1_28.inv_2  (    .in(\inv4_stage1_28.in ),    .out(\inv4_stage1_28.out )
  );
  inverter \inv4_stage1_28.inv_3  (    .in(\inv4_stage1_28.in ),    .out(\inv4_stage1_28.out )
  );
  inverter \inv4_stage1_29.inv_0  (    .in(\inv4_stage1_29.in ),    .out(\inv4_stage1_29.out )
  );
  inverter \inv4_stage1_29.inv_1  (    .in(\inv4_stage1_29.in ),    .out(\inv4_stage1_29.out )
  );
  inverter \inv4_stage1_29.inv_2  (    .in(\inv4_stage1_29.in ),    .out(\inv4_stage1_29.out )
  );
  inverter \inv4_stage1_29.inv_3  (    .in(\inv4_stage1_29.in ),    .out(\inv4_stage1_29.out )
  );
  inverter \inv4_stage1_3.inv_0  (    .in(\inv4_stage1_3.in ),    .out(\inv4_stage1_3.out )
  );
  inverter \inv4_stage1_3.inv_1  (    .in(\inv4_stage1_3.in ),    .out(\inv4_stage1_3.out )
  );
  inverter \inv4_stage1_3.inv_2  (    .in(\inv4_stage1_3.in ),    .out(\inv4_stage1_3.out )
  );
  inverter \inv4_stage1_3.inv_3  (    .in(\inv4_stage1_3.in ),    .out(\inv4_stage1_3.out )
  );
  inverter \inv4_stage1_30.inv_0  (    .in(\inv4_stage1_30.in ),    .out(\inv4_stage1_30.out )
  );
  inverter \inv4_stage1_30.inv_1  (    .in(\inv4_stage1_30.in ),    .out(\inv4_stage1_30.out )
  );
  inverter \inv4_stage1_30.inv_2  (    .in(\inv4_stage1_30.in ),    .out(\inv4_stage1_30.out )
  );
  inverter \inv4_stage1_30.inv_3  (    .in(\inv4_stage1_30.in ),    .out(\inv4_stage1_30.out )
  );
  inverter \inv4_stage1_31.inv_0  (    .in(\inv4_stage1_31.in ),    .out(\inv4_stage1_31.out )
  );
  inverter \inv4_stage1_31.inv_1  (    .in(\inv4_stage1_31.in ),    .out(\inv4_stage1_31.out )
  );
  inverter \inv4_stage1_31.inv_2  (    .in(\inv4_stage1_31.in ),    .out(\inv4_stage1_31.out )
  );
  inverter \inv4_stage1_31.inv_3  (    .in(\inv4_stage1_31.in ),    .out(\inv4_stage1_31.out )
  );
  inverter \inv4_stage1_32.inv_0  (    .in(\inv4_stage1_32.in ),    .out(\inv4_stage1_32.out )
  );
  inverter \inv4_stage1_32.inv_1  (    .in(\inv4_stage1_32.in ),    .out(\inv4_stage1_32.out )
  );
  inverter \inv4_stage1_32.inv_2  (    .in(\inv4_stage1_32.in ),    .out(\inv4_stage1_32.out )
  );
  inverter \inv4_stage1_32.inv_3  (    .in(\inv4_stage1_32.in ),    .out(\inv4_stage1_32.out )
  );
  inverter \inv4_stage1_33.inv_0  (    .in(\inv4_stage1_33.in ),    .out(\inv4_stage1_33.out )
  );
  inverter \inv4_stage1_33.inv_1  (    .in(\inv4_stage1_33.in ),    .out(\inv4_stage1_33.out )
  );
  inverter \inv4_stage1_33.inv_2  (    .in(\inv4_stage1_33.in ),    .out(\inv4_stage1_33.out )
  );
  inverter \inv4_stage1_33.inv_3  (    .in(\inv4_stage1_33.in ),    .out(\inv4_stage1_33.out )
  );
  inverter \inv4_stage1_34.inv_0  (    .in(\inv4_stage1_34.in ),    .out(\inv4_stage1_34.out )
  );
  inverter \inv4_stage1_34.inv_1  (    .in(\inv4_stage1_34.in ),    .out(\inv4_stage1_34.out )
  );
  inverter \inv4_stage1_34.inv_2  (    .in(\inv4_stage1_34.in ),    .out(\inv4_stage1_34.out )
  );
  inverter \inv4_stage1_34.inv_3  (    .in(\inv4_stage1_34.in ),    .out(\inv4_stage1_34.out )
  );
  inverter \inv4_stage1_35.inv_0  (    .in(\inv4_stage1_35.in ),    .out(\inv4_stage1_35.out )
  );
  inverter \inv4_stage1_35.inv_1  (    .in(\inv4_stage1_35.in ),    .out(\inv4_stage1_35.out )
  );
  inverter \inv4_stage1_35.inv_2  (    .in(\inv4_stage1_35.in ),    .out(\inv4_stage1_35.out )
  );
  inverter \inv4_stage1_35.inv_3  (    .in(\inv4_stage1_35.in ),    .out(\inv4_stage1_35.out )
  );
  inverter \inv4_stage1_36.inv_0  (    .in(\inv4_stage1_36.in ),    .out(\inv4_stage1_36.out )
  );
  inverter \inv4_stage1_36.inv_1  (    .in(\inv4_stage1_36.in ),    .out(\inv4_stage1_36.out )
  );
  inverter \inv4_stage1_36.inv_2  (    .in(\inv4_stage1_36.in ),    .out(\inv4_stage1_36.out )
  );
  inverter \inv4_stage1_36.inv_3  (    .in(\inv4_stage1_36.in ),    .out(\inv4_stage1_36.out )
  );
  inverter \inv4_stage1_37.inv_0  (    .in(\inv4_stage1_37.in ),    .out(\inv4_stage1_37.out )
  );
  inverter \inv4_stage1_37.inv_1  (    .in(\inv4_stage1_37.in ),    .out(\inv4_stage1_37.out )
  );
  inverter \inv4_stage1_37.inv_2  (    .in(\inv4_stage1_37.in ),    .out(\inv4_stage1_37.out )
  );
  inverter \inv4_stage1_37.inv_3  (    .in(\inv4_stage1_37.in ),    .out(\inv4_stage1_37.out )
  );
  inverter \inv4_stage1_38.inv_0  (    .in(\inv4_stage1_38.in ),    .out(\inv4_stage1_38.out )
  );
  inverter \inv4_stage1_38.inv_1  (    .in(\inv4_stage1_38.in ),    .out(\inv4_stage1_38.out )
  );
  inverter \inv4_stage1_38.inv_2  (    .in(\inv4_stage1_38.in ),    .out(\inv4_stage1_38.out )
  );
  inverter \inv4_stage1_38.inv_3  (    .in(\inv4_stage1_38.in ),    .out(\inv4_stage1_38.out )
  );
  inverter \inv4_stage1_39.inv_0  (    .in(\inv4_stage1_39.in ),    .out(\inv4_stage1_39.out )
  );
  inverter \inv4_stage1_39.inv_1  (    .in(\inv4_stage1_39.in ),    .out(\inv4_stage1_39.out )
  );
  inverter \inv4_stage1_39.inv_2  (    .in(\inv4_stage1_39.in ),    .out(\inv4_stage1_39.out )
  );
  inverter \inv4_stage1_39.inv_3  (    .in(\inv4_stage1_39.in ),    .out(\inv4_stage1_39.out )
  );
  inverter \inv4_stage1_4.inv_0  (    .in(\inv4_stage1_4.in ),    .out(\inv4_stage1_4.out )
  );
  inverter \inv4_stage1_4.inv_1  (    .in(\inv4_stage1_4.in ),    .out(\inv4_stage1_4.out )
  );
  inverter \inv4_stage1_4.inv_2  (    .in(\inv4_stage1_4.in ),    .out(\inv4_stage1_4.out )
  );
  inverter \inv4_stage1_4.inv_3  (    .in(\inv4_stage1_4.in ),    .out(\inv4_stage1_4.out )
  );
  inverter \inv4_stage1_40.inv_0  (    .in(\inv4_stage1_40.in ),    .out(\inv4_stage1_40.out )
  );
  inverter \inv4_stage1_40.inv_1  (    .in(\inv4_stage1_40.in ),    .out(\inv4_stage1_40.out )
  );
  inverter \inv4_stage1_40.inv_2  (    .in(\inv4_stage1_40.in ),    .out(\inv4_stage1_40.out )
  );
  inverter \inv4_stage1_40.inv_3  (    .in(\inv4_stage1_40.in ),    .out(\inv4_stage1_40.out )
  );
  inverter \inv4_stage1_41.inv_0  (    .in(\inv4_stage1_41.in ),    .out(\inv4_stage1_41.out )
  );
  inverter \inv4_stage1_41.inv_1  (    .in(\inv4_stage1_41.in ),    .out(\inv4_stage1_41.out )
  );
  inverter \inv4_stage1_41.inv_2  (    .in(\inv4_stage1_41.in ),    .out(\inv4_stage1_41.out )
  );
  inverter \inv4_stage1_41.inv_3  (    .in(\inv4_stage1_41.in ),    .out(\inv4_stage1_41.out )
  );
  inverter \inv4_stage1_42.inv_0  (    .in(\inv4_stage1_42.in ),    .out(\inv4_stage1_42.out )
  );
  inverter \inv4_stage1_42.inv_1  (    .in(\inv4_stage1_42.in ),    .out(\inv4_stage1_42.out )
  );
  inverter \inv4_stage1_42.inv_2  (    .in(\inv4_stage1_42.in ),    .out(\inv4_stage1_42.out )
  );
  inverter \inv4_stage1_42.inv_3  (    .in(\inv4_stage1_42.in ),    .out(\inv4_stage1_42.out )
  );
  inverter \inv4_stage1_43.inv_0  (    .in(\inv4_stage1_43.in ),    .out(\inv4_stage1_43.out )
  );
  inverter \inv4_stage1_43.inv_1  (    .in(\inv4_stage1_43.in ),    .out(\inv4_stage1_43.out )
  );
  inverter \inv4_stage1_43.inv_2  (    .in(\inv4_stage1_43.in ),    .out(\inv4_stage1_43.out )
  );
  inverter \inv4_stage1_43.inv_3  (    .in(\inv4_stage1_43.in ),    .out(\inv4_stage1_43.out )
  );
  inverter \inv4_stage1_44.inv_0  (    .in(\inv4_stage1_44.in ),    .out(\inv4_stage1_44.out )
  );
  inverter \inv4_stage1_44.inv_1  (    .in(\inv4_stage1_44.in ),    .out(\inv4_stage1_44.out )
  );
  inverter \inv4_stage1_44.inv_2  (    .in(\inv4_stage1_44.in ),    .out(\inv4_stage1_44.out )
  );
  inverter \inv4_stage1_44.inv_3  (    .in(\inv4_stage1_44.in ),    .out(\inv4_stage1_44.out )
  );
  inverter \inv4_stage1_45.inv_0  (    .in(\inv4_stage1_45.in ),    .out(\inv4_stage1_45.out )
  );
  inverter \inv4_stage1_45.inv_1  (    .in(\inv4_stage1_45.in ),    .out(\inv4_stage1_45.out )
  );
  inverter \inv4_stage1_45.inv_2  (    .in(\inv4_stage1_45.in ),    .out(\inv4_stage1_45.out )
  );
  inverter \inv4_stage1_45.inv_3  (    .in(\inv4_stage1_45.in ),    .out(\inv4_stage1_45.out )
  );
  inverter \inv4_stage1_46.inv_0  (    .in(\inv4_stage1_46.in ),    .out(\inv4_stage1_46.out )
  );
  inverter \inv4_stage1_46.inv_1  (    .in(\inv4_stage1_46.in ),    .out(\inv4_stage1_46.out )
  );
  inverter \inv4_stage1_46.inv_2  (    .in(\inv4_stage1_46.in ),    .out(\inv4_stage1_46.out )
  );
  inverter \inv4_stage1_46.inv_3  (    .in(\inv4_stage1_46.in ),    .out(\inv4_stage1_46.out )
  );
  inverter \inv4_stage1_47.inv_0  (    .in(\inv4_stage1_47.in ),    .out(\inv4_stage1_47.out )
  );
  inverter \inv4_stage1_47.inv_1  (    .in(\inv4_stage1_47.in ),    .out(\inv4_stage1_47.out )
  );
  inverter \inv4_stage1_47.inv_2  (    .in(\inv4_stage1_47.in ),    .out(\inv4_stage1_47.out )
  );
  inverter \inv4_stage1_47.inv_3  (    .in(\inv4_stage1_47.in ),    .out(\inv4_stage1_47.out )
  );
  inverter \inv4_stage1_48.inv_0  (    .in(\inv4_stage1_48.in ),    .out(\inv4_stage1_48.out )
  );
  inverter \inv4_stage1_48.inv_1  (    .in(\inv4_stage1_48.in ),    .out(\inv4_stage1_48.out )
  );
  inverter \inv4_stage1_48.inv_2  (    .in(\inv4_stage1_48.in ),    .out(\inv4_stage1_48.out )
  );
  inverter \inv4_stage1_48.inv_3  (    .in(\inv4_stage1_48.in ),    .out(\inv4_stage1_48.out )
  );
  inverter \inv4_stage1_49.inv_0  (    .in(\inv4_stage1_49.in ),    .out(\inv4_stage1_49.out )
  );
  inverter \inv4_stage1_49.inv_1  (    .in(\inv4_stage1_49.in ),    .out(\inv4_stage1_49.out )
  );
  inverter \inv4_stage1_49.inv_2  (    .in(\inv4_stage1_49.in ),    .out(\inv4_stage1_49.out )
  );
  inverter \inv4_stage1_49.inv_3  (    .in(\inv4_stage1_49.in ),    .out(\inv4_stage1_49.out )
  );
  inverter \inv4_stage1_5.inv_0  (    .in(\inv4_stage1_5.in ),    .out(\inv4_stage1_5.out )
  );
  inverter \inv4_stage1_5.inv_1  (    .in(\inv4_stage1_5.in ),    .out(\inv4_stage1_5.out )
  );
  inverter \inv4_stage1_5.inv_2  (    .in(\inv4_stage1_5.in ),    .out(\inv4_stage1_5.out )
  );
  inverter \inv4_stage1_5.inv_3  (    .in(\inv4_stage1_5.in ),    .out(\inv4_stage1_5.out )
  );
  inverter \inv4_stage1_50.inv_0  (    .in(\inv4_stage1_50.in ),    .out(\inv4_stage1_50.out )
  );
  inverter \inv4_stage1_50.inv_1  (    .in(\inv4_stage1_50.in ),    .out(\inv4_stage1_50.out )
  );
  inverter \inv4_stage1_50.inv_2  (    .in(\inv4_stage1_50.in ),    .out(\inv4_stage1_50.out )
  );
  inverter \inv4_stage1_50.inv_3  (    .in(\inv4_stage1_50.in ),    .out(\inv4_stage1_50.out )
  );
  inverter \inv4_stage1_51.inv_0  (    .in(\inv4_stage1_51.in ),    .out(\inv4_stage1_51.out )
  );
  inverter \inv4_stage1_51.inv_1  (    .in(\inv4_stage1_51.in ),    .out(\inv4_stage1_51.out )
  );
  inverter \inv4_stage1_51.inv_2  (    .in(\inv4_stage1_51.in ),    .out(\inv4_stage1_51.out )
  );
  inverter \inv4_stage1_51.inv_3  (    .in(\inv4_stage1_51.in ),    .out(\inv4_stage1_51.out )
  );
  inverter \inv4_stage1_52.inv_0  (    .in(\inv4_stage1_52.in ),    .out(\inv4_stage1_52.out )
  );
  inverter \inv4_stage1_52.inv_1  (    .in(\inv4_stage1_52.in ),    .out(\inv4_stage1_52.out )
  );
  inverter \inv4_stage1_52.inv_2  (    .in(\inv4_stage1_52.in ),    .out(\inv4_stage1_52.out )
  );
  inverter \inv4_stage1_52.inv_3  (    .in(\inv4_stage1_52.in ),    .out(\inv4_stage1_52.out )
  );
  inverter \inv4_stage1_53.inv_0  (    .in(\inv4_stage1_53.in ),    .out(\inv4_stage1_53.out )
  );
  inverter \inv4_stage1_53.inv_1  (    .in(\inv4_stage1_53.in ),    .out(\inv4_stage1_53.out )
  );
  inverter \inv4_stage1_53.inv_2  (    .in(\inv4_stage1_53.in ),    .out(\inv4_stage1_53.out )
  );
  inverter \inv4_stage1_53.inv_3  (    .in(\inv4_stage1_53.in ),    .out(\inv4_stage1_53.out )
  );
  inverter \inv4_stage1_54.inv_0  (    .in(\inv4_stage1_54.in ),    .out(\inv4_stage1_54.out )
  );
  inverter \inv4_stage1_54.inv_1  (    .in(\inv4_stage1_54.in ),    .out(\inv4_stage1_54.out )
  );
  inverter \inv4_stage1_54.inv_2  (    .in(\inv4_stage1_54.in ),    .out(\inv4_stage1_54.out )
  );
  inverter \inv4_stage1_54.inv_3  (    .in(\inv4_stage1_54.in ),    .out(\inv4_stage1_54.out )
  );
  inverter \inv4_stage1_55.inv_0  (    .in(\inv4_stage1_55.in ),    .out(\inv4_stage1_55.out )
  );
  inverter \inv4_stage1_55.inv_1  (    .in(\inv4_stage1_55.in ),    .out(\inv4_stage1_55.out )
  );
  inverter \inv4_stage1_55.inv_2  (    .in(\inv4_stage1_55.in ),    .out(\inv4_stage1_55.out )
  );
  inverter \inv4_stage1_55.inv_3  (    .in(\inv4_stage1_55.in ),    .out(\inv4_stage1_55.out )
  );
  inverter \inv4_stage1_56.inv_0  (    .in(\inv4_stage1_56.in ),    .out(\inv4_stage1_56.out )
  );
  inverter \inv4_stage1_56.inv_1  (    .in(\inv4_stage1_56.in ),    .out(\inv4_stage1_56.out )
  );
  inverter \inv4_stage1_56.inv_2  (    .in(\inv4_stage1_56.in ),    .out(\inv4_stage1_56.out )
  );
  inverter \inv4_stage1_56.inv_3  (    .in(\inv4_stage1_56.in ),    .out(\inv4_stage1_56.out )
  );
  inverter \inv4_stage1_57.inv_0  (    .in(\inv4_stage1_57.in ),    .out(\inv4_stage1_57.out )
  );
  inverter \inv4_stage1_57.inv_1  (    .in(\inv4_stage1_57.in ),    .out(\inv4_stage1_57.out )
  );
  inverter \inv4_stage1_57.inv_2  (    .in(\inv4_stage1_57.in ),    .out(\inv4_stage1_57.out )
  );
  inverter \inv4_stage1_57.inv_3  (    .in(\inv4_stage1_57.in ),    .out(\inv4_stage1_57.out )
  );
  inverter \inv4_stage1_58.inv_0  (    .in(\inv4_stage1_58.in ),    .out(\inv4_stage1_58.out )
  );
  inverter \inv4_stage1_58.inv_1  (    .in(\inv4_stage1_58.in ),    .out(\inv4_stage1_58.out )
  );
  inverter \inv4_stage1_58.inv_2  (    .in(\inv4_stage1_58.in ),    .out(\inv4_stage1_58.out )
  );
  inverter \inv4_stage1_58.inv_3  (    .in(\inv4_stage1_58.in ),    .out(\inv4_stage1_58.out )
  );
  inverter \inv4_stage1_59.inv_0  (    .in(\inv4_stage1_59.in ),    .out(\inv4_stage1_59.out )
  );
  inverter \inv4_stage1_59.inv_1  (    .in(\inv4_stage1_59.in ),    .out(\inv4_stage1_59.out )
  );
  inverter \inv4_stage1_59.inv_2  (    .in(\inv4_stage1_59.in ),    .out(\inv4_stage1_59.out )
  );
  inverter \inv4_stage1_59.inv_3  (    .in(\inv4_stage1_59.in ),    .out(\inv4_stage1_59.out )
  );
  inverter \inv4_stage1_6.inv_0  (    .in(\inv4_stage1_6.in ),    .out(\inv4_stage1_6.out )
  );
  inverter \inv4_stage1_6.inv_1  (    .in(\inv4_stage1_6.in ),    .out(\inv4_stage1_6.out )
  );
  inverter \inv4_stage1_6.inv_2  (    .in(\inv4_stage1_6.in ),    .out(\inv4_stage1_6.out )
  );
  inverter \inv4_stage1_6.inv_3  (    .in(\inv4_stage1_6.in ),    .out(\inv4_stage1_6.out )
  );
  inverter \inv4_stage1_60.inv_0  (    .in(\inv4_stage1_60.in ),    .out(\inv4_stage1_60.out )
  );
  inverter \inv4_stage1_60.inv_1  (    .in(\inv4_stage1_60.in ),    .out(\inv4_stage1_60.out )
  );
  inverter \inv4_stage1_60.inv_2  (    .in(\inv4_stage1_60.in ),    .out(\inv4_stage1_60.out )
  );
  inverter \inv4_stage1_60.inv_3  (    .in(\inv4_stage1_60.in ),    .out(\inv4_stage1_60.out )
  );
  inverter \inv4_stage1_61.inv_0  (    .in(\inv4_stage1_61.in ),    .out(\inv4_stage1_61.out )
  );
  inverter \inv4_stage1_61.inv_1  (    .in(\inv4_stage1_61.in ),    .out(\inv4_stage1_61.out )
  );
  inverter \inv4_stage1_61.inv_2  (    .in(\inv4_stage1_61.in ),    .out(\inv4_stage1_61.out )
  );
  inverter \inv4_stage1_61.inv_3  (    .in(\inv4_stage1_61.in ),    .out(\inv4_stage1_61.out )
  );
  inverter \inv4_stage1_62.inv_0  (    .in(\inv4_stage1_62.in ),    .out(\inv4_stage1_62.out )
  );
  inverter \inv4_stage1_62.inv_1  (    .in(\inv4_stage1_62.in ),    .out(\inv4_stage1_62.out )
  );
  inverter \inv4_stage1_62.inv_2  (    .in(\inv4_stage1_62.in ),    .out(\inv4_stage1_62.out )
  );
  inverter \inv4_stage1_62.inv_3  (    .in(\inv4_stage1_62.in ),    .out(\inv4_stage1_62.out )
  );
  inverter \inv4_stage1_63.inv_0  (    .in(\inv4_stage1_63.in ),    .out(\inv4_stage1_63.out )
  );
  inverter \inv4_stage1_63.inv_1  (    .in(\inv4_stage1_63.in ),    .out(\inv4_stage1_63.out )
  );
  inverter \inv4_stage1_63.inv_2  (    .in(\inv4_stage1_63.in ),    .out(\inv4_stage1_63.out )
  );
  inverter \inv4_stage1_63.inv_3  (    .in(\inv4_stage1_63.in ),    .out(\inv4_stage1_63.out )
  );
  inverter \inv4_stage1_7.inv_0  (    .in(\inv4_stage1_7.in ),    .out(\inv4_stage1_7.out )
  );
  inverter \inv4_stage1_7.inv_1  (    .in(\inv4_stage1_7.in ),    .out(\inv4_stage1_7.out )
  );
  inverter \inv4_stage1_7.inv_2  (    .in(\inv4_stage1_7.in ),    .out(\inv4_stage1_7.out )
  );
  inverter \inv4_stage1_7.inv_3  (    .in(\inv4_stage1_7.in ),    .out(\inv4_stage1_7.out )
  );
  inverter \inv4_stage1_8.inv_0  (    .in(\inv4_stage1_8.in ),    .out(\inv4_stage1_8.out )
  );
  inverter \inv4_stage1_8.inv_1  (    .in(\inv4_stage1_8.in ),    .out(\inv4_stage1_8.out )
  );
  inverter \inv4_stage1_8.inv_2  (    .in(\inv4_stage1_8.in ),    .out(\inv4_stage1_8.out )
  );
  inverter \inv4_stage1_8.inv_3  (    .in(\inv4_stage1_8.in ),    .out(\inv4_stage1_8.out )
  );
  inverter \inv4_stage1_9.inv_0  (    .in(\inv4_stage1_9.in ),    .out(\inv4_stage1_9.out )
  );
  inverter \inv4_stage1_9.inv_1  (    .in(\inv4_stage1_9.in ),    .out(\inv4_stage1_9.out )
  );
  inverter \inv4_stage1_9.inv_2  (    .in(\inv4_stage1_9.in ),    .out(\inv4_stage1_9.out )
  );
  inverter \inv4_stage1_9.inv_3  (    .in(\inv4_stage1_9.in ),    .out(\inv4_stage1_9.out )
  );
  inverter inv_stage0_0 (    .in(\in<0> ),    .out(\inv4_stage1_0.in )
  );
  inverter inv_stage0_1 (    .in(\in<1> ),    .out(\inv4_stage1_1.in )
  );
  inverter inv_stage0_10 (    .in(\in<10> ),    .out(\inv4_stage1_10.in )
  );
  inverter inv_stage0_11 (    .in(\in<11> ),    .out(\inv4_stage1_11.in )
  );
  inverter inv_stage0_12 (    .in(\in<12> ),    .out(\inv4_stage1_12.in )
  );
  inverter inv_stage0_13 (    .in(\in<13> ),    .out(\inv4_stage1_13.in )
  );
  inverter inv_stage0_14 (    .in(\in<14> ),    .out(\inv4_stage1_14.in )
  );
  inverter inv_stage0_15 (    .in(\in<15> ),    .out(\inv4_stage1_15.in )
  );
  inverter inv_stage0_16 (    .in(\in<16> ),    .out(\inv4_stage1_16.in )
  );
  inverter inv_stage0_17 (    .in(\in<17> ),    .out(\inv4_stage1_17.in )
  );
  inverter inv_stage0_18 (    .in(\in<18> ),    .out(\inv4_stage1_18.in )
  );
  inverter inv_stage0_19 (    .in(\in<19> ),    .out(\inv4_stage1_19.in )
  );
  inverter inv_stage0_2 (    .in(\in<2> ),    .out(\inv4_stage1_2.in )
  );
  inverter inv_stage0_20 (    .in(\in<20> ),    .out(\inv4_stage1_20.in )
  );
  inverter inv_stage0_21 (    .in(\in<21> ),    .out(\inv4_stage1_21.in )
  );
  inverter inv_stage0_22 (    .in(\in<22> ),    .out(\inv4_stage1_22.in )
  );
  inverter inv_stage0_23 (    .in(\in<23> ),    .out(\inv4_stage1_23.in )
  );
  inverter inv_stage0_24 (    .in(\in<24> ),    .out(\inv4_stage1_24.in )
  );
  inverter inv_stage0_25 (    .in(\in<25> ),    .out(\inv4_stage1_25.in )
  );
  inverter inv_stage0_26 (    .in(\in<26> ),    .out(\inv4_stage1_26.in )
  );
  inverter inv_stage0_27 (    .in(\in<27> ),    .out(\inv4_stage1_27.in )
  );
  inverter inv_stage0_28 (    .in(\in<28> ),    .out(\inv4_stage1_28.in )
  );
  inverter inv_stage0_29 (    .in(\in<29> ),    .out(\inv4_stage1_29.in )
  );
  inverter inv_stage0_3 (    .in(\in<3> ),    .out(\inv4_stage1_3.in )
  );
  inverter inv_stage0_30 (    .in(\in<30> ),    .out(\inv4_stage1_30.in )
  );
  inverter inv_stage0_31 (    .in(\in<31> ),    .out(\inv4_stage1_31.in )
  );
  inverter inv_stage0_32 (    .in(\in<32> ),    .out(\inv4_stage1_32.in )
  );
  inverter inv_stage0_33 (    .in(\in<33> ),    .out(\inv4_stage1_33.in )
  );
  inverter inv_stage0_34 (    .in(\in<34> ),    .out(\inv4_stage1_34.in )
  );
  inverter inv_stage0_35 (    .in(\in<35> ),    .out(\inv4_stage1_35.in )
  );
  inverter inv_stage0_36 (    .in(\in<36> ),    .out(\inv4_stage1_36.in )
  );
  inverter inv_stage0_37 (    .in(\in<37> ),    .out(\inv4_stage1_37.in )
  );
  inverter inv_stage0_38 (    .in(\in<38> ),    .out(\inv4_stage1_38.in )
  );
  inverter inv_stage0_39 (    .in(\in<39> ),    .out(\inv4_stage1_39.in )
  );
  inverter inv_stage0_4 (    .in(\in<4> ),    .out(\inv4_stage1_4.in )
  );
  inverter inv_stage0_40 (    .in(\in<40> ),    .out(\inv4_stage1_40.in )
  );
  inverter inv_stage0_41 (    .in(\in<41> ),    .out(\inv4_stage1_41.in )
  );
  inverter inv_stage0_42 (    .in(\in<42> ),    .out(\inv4_stage1_42.in )
  );
  inverter inv_stage0_43 (    .in(\in<43> ),    .out(\inv4_stage1_43.in )
  );
  inverter inv_stage0_44 (    .in(\in<44> ),    .out(\inv4_stage1_44.in )
  );
  inverter inv_stage0_45 (    .in(\in<45> ),    .out(\inv4_stage1_45.in )
  );
  inverter inv_stage0_46 (    .in(\in<46> ),    .out(\inv4_stage1_46.in )
  );
  inverter inv_stage0_47 (    .in(\in<47> ),    .out(\inv4_stage1_47.in )
  );
  inverter inv_stage0_48 (    .in(\in<48> ),    .out(\inv4_stage1_48.in )
  );
  inverter inv_stage0_49 (    .in(\in<49> ),    .out(\inv4_stage1_49.in )
  );
  inverter inv_stage0_5 (    .in(\in<5> ),    .out(\inv4_stage1_5.in )
  );
  inverter inv_stage0_50 (    .in(\in<50> ),    .out(\inv4_stage1_50.in )
  );
  inverter inv_stage0_51 (    .in(\in<51> ),    .out(\inv4_stage1_51.in )
  );
  inverter inv_stage0_52 (    .in(\in<52> ),    .out(\inv4_stage1_52.in )
  );
  inverter inv_stage0_53 (    .in(\in<53> ),    .out(\inv4_stage1_53.in )
  );
  inverter inv_stage0_54 (    .in(\in<54> ),    .out(\inv4_stage1_54.in )
  );
  inverter inv_stage0_55 (    .in(\in<55> ),    .out(\inv4_stage1_55.in )
  );
  inverter inv_stage0_56 (    .in(\in<56> ),    .out(\inv4_stage1_56.in )
  );
  inverter inv_stage0_57 (    .in(\in<57> ),    .out(\inv4_stage1_57.in )
  );
  inverter inv_stage0_58 (    .in(\in<58> ),    .out(\inv4_stage1_58.in )
  );
  inverter inv_stage0_59 (    .in(\in<59> ),    .out(\inv4_stage1_59.in )
  );
  inverter inv_stage0_6 (    .in(\in<6> ),    .out(\inv4_stage1_6.in )
  );
  inverter inv_stage0_60 (    .in(\in<60> ),    .out(\inv4_stage1_60.in )
  );
  inverter inv_stage0_61 (    .in(\in<61> ),    .out(\inv4_stage1_61.in )
  );
  inverter inv_stage0_62 (    .in(\in<62> ),    .out(\inv4_stage1_62.in )
  );
  inverter inv_stage0_63 (    .in(\in<63> ),    .out(\inv4_stage1_63.in )
  );
  inverter inv_stage0_7 (    .in(\in<7> ),    .out(\inv4_stage1_7.in )
  );
  inverter inv_stage0_8 (    .in(\in<8> ),    .out(\inv4_stage1_8.in )
  );
  inverter inv_stage0_9 (    .in(\in<9> ),    .out(\inv4_stage1_9.in )
  );
  assign \out_b<63>  = \inv4_stage1_63.in ;
  assign \out_b<62>  = \inv4_stage1_62.in ;
  assign \out_b<61>  = \inv4_stage1_61.in ;
  assign \out_b<60>  = \inv4_stage1_60.in ;
  assign \out_b<59>  = \inv4_stage1_59.in ;
  assign \out_b<58>  = \inv4_stage1_58.in ;
  assign \out_b<57>  = \inv4_stage1_57.in ;
  assign \out_b<56>  = \inv4_stage1_56.in ;
  assign \out_b<55>  = \inv4_stage1_55.in ;
  assign \out_b<54>  = \inv4_stage1_54.in ;
  assign \out_b<53>  = \inv4_stage1_53.in ;
  assign \out_b<52>  = \inv4_stage1_52.in ;
  assign \out_b<51>  = \inv4_stage1_51.in ;
  assign \out_b<50>  = \inv4_stage1_50.in ;
  assign \out_b<49>  = \inv4_stage1_49.in ;
  assign \out_b<48>  = \inv4_stage1_48.in ;
  assign \out_b<47>  = \inv4_stage1_47.in ;
  assign \out_b<46>  = \inv4_stage1_46.in ;
  assign \out_b<45>  = \inv4_stage1_45.in ;
  assign \out_b<44>  = \inv4_stage1_44.in ;
  assign \out_b<43>  = \inv4_stage1_43.in ;
  assign \out_b<42>  = \inv4_stage1_42.in ;
  assign \out_b<41>  = \inv4_stage1_41.in ;
  assign \out_b<40>  = \inv4_stage1_40.in ;
  assign \out_b<39>  = \inv4_stage1_39.in ;
  assign \out_b<38>  = \inv4_stage1_38.in ;
  assign \out_b<37>  = \inv4_stage1_37.in ;
  assign \out_b<36>  = \inv4_stage1_36.in ;
  assign \out_b<35>  = \inv4_stage1_35.in ;
  assign \out_b<34>  = \inv4_stage1_34.in ;
  assign \out_b<33>  = \inv4_stage1_33.in ;
  assign \out_b<32>  = \inv4_stage1_32.in ;
  assign \out_b<31>  = \inv4_stage1_31.in ;
  assign \out_b<30>  = \inv4_stage1_30.in ;
  assign \out_b<29>  = \inv4_stage1_29.in ;
  assign \out_b<28>  = \inv4_stage1_28.in ;
  assign \out_b<27>  = \inv4_stage1_27.in ;
  assign \out_b<26>  = \inv4_stage1_26.in ;
  assign \out_b<25>  = \inv4_stage1_25.in ;
  assign \out_b<24>  = \inv4_stage1_24.in ;
  assign \out_b<23>  = \inv4_stage1_23.in ;
  assign \out_b<22>  = \inv4_stage1_22.in ;
  assign \out_b<21>  = \inv4_stage1_21.in ;
  assign \out_b<20>  = \inv4_stage1_20.in ;
  assign \out_b<19>  = \inv4_stage1_19.in ;
  assign \out_b<18>  = \inv4_stage1_18.in ;
  assign \out_b<17>  = \inv4_stage1_17.in ;
  assign \out_b<16>  = \inv4_stage1_16.in ;
  assign \out_b<15>  = \inv4_stage1_15.in ;
  assign \out_b<14>  = \inv4_stage1_14.in ;
  assign \out_b<13>  = \inv4_stage1_13.in ;
  assign \out_b<12>  = \inv4_stage1_12.in ;
  assign \out_b<11>  = \inv4_stage1_11.in ;
  assign \out_b<10>  = \inv4_stage1_10.in ;
  assign \out_b<9>  = \inv4_stage1_9.in ;
  assign \out_b<8>  = \inv4_stage1_8.in ;
  assign \out_b<7>  = \inv4_stage1_7.in ;
  assign \out_b<6>  = \inv4_stage1_6.in ;
  assign \out_b<5>  = \inv4_stage1_5.in ;
  assign \out_b<4>  = \inv4_stage1_4.in ;
  assign \out_b<3>  = \inv4_stage1_3.in ;
  assign \out_b<2>  = \inv4_stage1_2.in ;
  assign \out_b<1>  = \inv4_stage1_1.in ;
  assign \out_b<0>  = \inv4_stage1_0.in ;
  assign \out<63>  = \inv4_stage1_63.out ;
  assign \out<62>  = \inv4_stage1_62.out ;
  assign \out<61>  = \inv4_stage1_61.out ;
  assign \out<60>  = \inv4_stage1_60.out ;
  assign \out<59>  = \inv4_stage1_59.out ;
  assign \out<58>  = \inv4_stage1_58.out ;
  assign \out<57>  = \inv4_stage1_57.out ;
  assign \out<56>  = \inv4_stage1_56.out ;
  assign \out<55>  = \inv4_stage1_55.out ;
  assign \out<54>  = \inv4_stage1_54.out ;
  assign \out<53>  = \inv4_stage1_53.out ;
  assign \out<52>  = \inv4_stage1_52.out ;
  assign \out<51>  = \inv4_stage1_51.out ;
  assign \out<50>  = \inv4_stage1_50.out ;
  assign \out<49>  = \inv4_stage1_49.out ;
  assign \out<48>  = \inv4_stage1_48.out ;
  assign \out<47>  = \inv4_stage1_47.out ;
  assign \out<46>  = \inv4_stage1_46.out ;
  assign \out<45>  = \inv4_stage1_45.out ;
  assign \out<44>  = \inv4_stage1_44.out ;
  assign \out<43>  = \inv4_stage1_43.out ;
  assign \out<42>  = \inv4_stage1_42.out ;
  assign \out<41>  = \inv4_stage1_41.out ;
  assign \out<40>  = \inv4_stage1_40.out ;
  assign \out<39>  = \inv4_stage1_39.out ;
  assign \out<38>  = \inv4_stage1_38.out ;
  assign \out<37>  = \inv4_stage1_37.out ;
  assign \out<36>  = \inv4_stage1_36.out ;
  assign \out<35>  = \inv4_stage1_35.out ;
  assign \out<34>  = \inv4_stage1_34.out ;
  assign \out<33>  = \inv4_stage1_33.out ;
  assign \out<32>  = \inv4_stage1_32.out ;
  assign \out<31>  = \inv4_stage1_31.out ;
  assign \out<30>  = \inv4_stage1_30.out ;
  assign \out<29>  = \inv4_stage1_29.out ;
  assign \out<28>  = \inv4_stage1_28.out ;
  assign \out<27>  = \inv4_stage1_27.out ;
  assign \out<26>  = \inv4_stage1_26.out ;
  assign \out<25>  = \inv4_stage1_25.out ;
  assign \out<24>  = \inv4_stage1_24.out ;
  assign \out<23>  = \inv4_stage1_23.out ;
  assign \out<22>  = \inv4_stage1_22.out ;
  assign \out<21>  = \inv4_stage1_21.out ;
  assign \out<20>  = \inv4_stage1_20.out ;
  assign \out<19>  = \inv4_stage1_19.out ;
  assign \out<18>  = \inv4_stage1_18.out ;
  assign \out<17>  = \inv4_stage1_17.out ;
  assign \out<16>  = \inv4_stage1_16.out ;
  assign \out<15>  = \inv4_stage1_15.out ;
  assign \out<14>  = \inv4_stage1_14.out ;
  assign \out<13>  = \inv4_stage1_13.out ;
  assign \out<12>  = \inv4_stage1_12.out ;
  assign \out<11>  = \inv4_stage1_11.out ;
  assign \out<10>  = \inv4_stage1_10.out ;
  assign \out<9>  = \inv4_stage1_9.out ;
  assign \out<8>  = \inv4_stage1_8.out ;
  assign \out<7>  = \inv4_stage1_7.out ;
  assign \out<6>  = \inv4_stage1_6.out ;
  assign \out<5>  = \inv4_stage1_5.out ;
  assign \out<4>  = \inv4_stage1_4.out ;
  assign \out<3>  = \inv4_stage1_3.out ;
  assign \out<2>  = \inv4_stage1_2.out ;
  assign \out<1>  = \inv4_stage1_1.out ;
  assign \out<0>  = \inv4_stage1_0.out ;
endmodule
