
module adder_tree_4bit_to_10bit(sign_weight, \in_0<0> , \in_0<1> , \in_0<2> , \in_0<3> , \in_1<0> , \in_1<1> , \in_1<2> , \in_1<3> , \in_2<0> , \in_2<1> , \in_2<2> , \in_2<3> , \in_3<0> , \in_3<1> , \in_3<2> , \in_3<3> , \in_4<0> , \in_4<1> , \in_4<2> , \in_4<3> , \in_5<0> , \in_5<1> , \in_5<2> , \in_5<3> , \in_6<0> , \in_6<1> , \in_6<2> , \in_6<3> , \in_7<0> , \in_7<1> , \in_7<2> , \in_7<3> , \in_8<0> , \in_8<1> , \in_8<2> , \in_8<3> , \in_9<0> , \in_9<1> , \in_9<2> , \in_9<3> , \in_10<0> , \in_10<1> , \in_10<2> , \in_10<3> , \in_11<0> , \in_11<1> , \in_11<2> , \in_11<3> , \in_12<0> , \in_12<1> , \in_12<2> , \in_12<3> , \in_13<0> , \in_13<1> , \in_13<2> , \in_13<3> , \in_14<0> , \in_14<1> , \in_14<2> , \in_14<3> , \in_15<0> , \in_15<1> , \in_15<2> , \in_15<3> , \in_16<0> , \in_16<1> , \in_16<2> , \in_16<3> , \in_17<0> , \in_17<1> , \in_17<2> , \in_17<3> , \in_18<0> , \in_18<1> , \in_18<2> , \in_18<3> , \in_19<0> , \in_19<1> , \in_19<2> , \in_19<3> , \in_20<0> , \in_20<1> , \in_20<2> , \in_20<3> , \in_21<0> , \in_21<1> , \in_21<2> , \in_21<3> , \in_22<0> , \in_22<1> , \in_22<2> , \in_22<3> , \in_23<0> , \in_23<1> , \in_23<2> , \in_23<3> , \in_24<0> , \in_24<1> , \in_24<2> , \in_24<3> , \in_25<0> , \in_25<1> , \in_25<2> , \in_25<3> , \in_26<0> , \in_26<1> , \in_26<2> , \in_26<3> , \in_27<0> , \in_27<1> , \in_27<2> , \in_27<3> , \in_28<0> , \in_28<1> , \in_28<2> , \in_28<3> , \in_29<0> , \in_29<1> , \in_29<2> , \in_29<3> , \in_30<0> , \in_30<1> , \in_30<2> , \in_30<3> , \in_31<0> , \in_31<1> , \in_31<2> , \in_31<3> , \in_32<0> , \in_32<1> , \in_32<2> , \in_32<3> , \in_33<0> , \in_33<1> , \in_33<2> , \in_33<3> , \in_34<0> , \in_34<1> , \in_34<2> , \in_34<3> , \in_35<0> , \in_35<1> , \in_35<2> , \in_35<3> , \in_36<0> , \in_36<1> , \in_36<2> , \in_36<3> , \in_37<0> , \in_37<1> , \in_37<2> , \in_37<3> , \in_38<0> , \in_38<1> , \in_38<2> , \in_38<3> , \in_39<0> , \in_39<1> , \in_39<2> , \in_39<3> , \in_40<0> , \in_40<1> , \in_40<2> , \in_40<3> , \in_41<0> , \in_41<1> , \in_41<2> , \in_41<3> , \in_42<0> , \in_42<1> , \in_42<2> , \in_42<3> , \in_43<0> , \in_43<1> , \in_43<2> , \in_43<3> , \in_44<0> , \in_44<1> , \in_44<2> , \in_44<3> , \in_45<0> , \in_45<1> , \in_45<2> , \in_45<3> , \in_46<0> , \in_46<1> , \in_46<2> , \in_46<3> , \in_47<0> , \in_47<1> , \in_47<2> , \in_47<3> , \in_48<0> , \in_48<1> , \in_48<2> , \in_48<3> , \in_49<0> , \in_49<1> , \in_49<2> , \in_49<3> , \in_50<0> , \in_50<1> , \in_50<2> , \in_50<3> , \in_51<0> , \in_51<1> , \in_51<2> , \in_51<3> , \in_52<0> , \in_52<1> , \in_52<2> , \in_52<3> , \in_53<0> , \in_53<1> , \in_53<2> , \in_53<3> , \in_54<0> , \in_54<1> , \in_54<2> , \in_54<3> , \in_55<0> , \in_55<1> , \in_55<2> , \in_55<3> , \in_56<0> , \in_56<1> , \in_56<2> , \in_56<3> , \in_57<0> , \in_57<1> , \in_57<2> , \in_57<3> , \in_58<0> , \in_58<1> , \in_58<2> , \in_58<3> , \in_59<0> , \in_59<1> , \in_59<2> , \in_59<3> , \in_60<0> , \in_60<1> , \in_60<2> , \in_60<3> , \in_61<0> , \in_61<1> , \in_61<2> , \in_61<3> , \in_62<0> , \in_62<1> , \in_62<2> , \in_62<3> , \in_63<0> , \in_63<1> , \in_63<2> , \in_63<3> , \out<0> , \out<1> , \out<2> , \out<3> , \out<4> , \out<5> , \out<6> , \out<7> , \out<8> , \out<9> );
  wire \adder_4bit_0.a<0> ;
  wire \adder_4bit_0.a<1> ;
  wire \adder_4bit_0.a<2> ;
  wire \adder_4bit_0.a<3> ;
  wire \adder_4bit_0.b<0> ;
  wire \adder_4bit_0.b<1> ;
  wire \adder_4bit_0.b<2> ;
  wire \adder_4bit_0.b<3> ;
  wire \adder_4bit_0.c<0> ;
  wire \adder_4bit_0.c<1> ;
  wire \adder_4bit_0.c<2> ;
  wire \adder_4bit_0.c<3> ;
  wire \adder_4bit_0.s<0> ;
  wire \adder_4bit_0.s<1> ;
  wire \adder_4bit_0.s<2> ;
  wire \adder_4bit_0.s<3> ;
  wire \adder_4bit_0.s<4> ;
  wire \adder_4bit_0.sign ;
  wire \adder_4bit_1.a<0> ;
  wire \adder_4bit_1.a<1> ;
  wire \adder_4bit_1.a<2> ;
  wire \adder_4bit_1.a<3> ;
  wire \adder_4bit_1.b<0> ;
  wire \adder_4bit_1.b<1> ;
  wire \adder_4bit_1.b<2> ;
  wire \adder_4bit_1.b<3> ;
  wire \adder_4bit_1.c<0> ;
  wire \adder_4bit_1.c<1> ;
  wire \adder_4bit_1.c<2> ;
  wire \adder_4bit_1.c<3> ;
  wire \adder_4bit_1.s<0> ;
  wire \adder_4bit_1.s<1> ;
  wire \adder_4bit_1.s<2> ;
  wire \adder_4bit_1.s<3> ;
  wire \adder_4bit_1.s<4> ;
  wire \adder_4bit_1.sign ;
  wire \adder_4bit_10.a<0> ;
  wire \adder_4bit_10.a<1> ;
  wire \adder_4bit_10.a<2> ;
  wire \adder_4bit_10.a<3> ;
  wire \adder_4bit_10.b<0> ;
  wire \adder_4bit_10.b<1> ;
  wire \adder_4bit_10.b<2> ;
  wire \adder_4bit_10.b<3> ;
  wire \adder_4bit_10.c<0> ;
  wire \adder_4bit_10.c<1> ;
  wire \adder_4bit_10.c<2> ;
  wire \adder_4bit_10.c<3> ;
  wire \adder_4bit_10.s<0> ;
  wire \adder_4bit_10.s<1> ;
  wire \adder_4bit_10.s<2> ;
  wire \adder_4bit_10.s<3> ;
  wire \adder_4bit_10.s<4> ;
  wire \adder_4bit_10.sign ;
  wire \adder_4bit_11.a<0> ;
  wire \adder_4bit_11.a<1> ;
  wire \adder_4bit_11.a<2> ;
  wire \adder_4bit_11.a<3> ;
  wire \adder_4bit_11.b<0> ;
  wire \adder_4bit_11.b<1> ;
  wire \adder_4bit_11.b<2> ;
  wire \adder_4bit_11.b<3> ;
  wire \adder_4bit_11.c<0> ;
  wire \adder_4bit_11.c<1> ;
  wire \adder_4bit_11.c<2> ;
  wire \adder_4bit_11.c<3> ;
  wire \adder_4bit_11.s<0> ;
  wire \adder_4bit_11.s<1> ;
  wire \adder_4bit_11.s<2> ;
  wire \adder_4bit_11.s<3> ;
  wire \adder_4bit_11.s<4> ;
  wire \adder_4bit_11.sign ;
  wire \adder_4bit_12.a<0> ;
  wire \adder_4bit_12.a<1> ;
  wire \adder_4bit_12.a<2> ;
  wire \adder_4bit_12.a<3> ;
  wire \adder_4bit_12.b<0> ;
  wire \adder_4bit_12.b<1> ;
  wire \adder_4bit_12.b<2> ;
  wire \adder_4bit_12.b<3> ;
  wire \adder_4bit_12.c<0> ;
  wire \adder_4bit_12.c<1> ;
  wire \adder_4bit_12.c<2> ;
  wire \adder_4bit_12.c<3> ;
  wire \adder_4bit_12.s<0> ;
  wire \adder_4bit_12.s<1> ;
  wire \adder_4bit_12.s<2> ;
  wire \adder_4bit_12.s<3> ;
  wire \adder_4bit_12.s<4> ;
  wire \adder_4bit_12.sign ;
  wire \adder_4bit_13.a<0> ;
  wire \adder_4bit_13.a<1> ;
  wire \adder_4bit_13.a<2> ;
  wire \adder_4bit_13.a<3> ;
  wire \adder_4bit_13.b<0> ;
  wire \adder_4bit_13.b<1> ;
  wire \adder_4bit_13.b<2> ;
  wire \adder_4bit_13.b<3> ;
  wire \adder_4bit_13.c<0> ;
  wire \adder_4bit_13.c<1> ;
  wire \adder_4bit_13.c<2> ;
  wire \adder_4bit_13.c<3> ;
  wire \adder_4bit_13.s<0> ;
  wire \adder_4bit_13.s<1> ;
  wire \adder_4bit_13.s<2> ;
  wire \adder_4bit_13.s<3> ;
  wire \adder_4bit_13.s<4> ;
  wire \adder_4bit_13.sign ;
  wire \adder_4bit_14.a<0> ;
  wire \adder_4bit_14.a<1> ;
  wire \adder_4bit_14.a<2> ;
  wire \adder_4bit_14.a<3> ;
  wire \adder_4bit_14.b<0> ;
  wire \adder_4bit_14.b<1> ;
  wire \adder_4bit_14.b<2> ;
  wire \adder_4bit_14.b<3> ;
  wire \adder_4bit_14.c<0> ;
  wire \adder_4bit_14.c<1> ;
  wire \adder_4bit_14.c<2> ;
  wire \adder_4bit_14.c<3> ;
  wire \adder_4bit_14.s<0> ;
  wire \adder_4bit_14.s<1> ;
  wire \adder_4bit_14.s<2> ;
  wire \adder_4bit_14.s<3> ;
  wire \adder_4bit_14.s<4> ;
  wire \adder_4bit_14.sign ;
  wire \adder_4bit_15.a<0> ;
  wire \adder_4bit_15.a<1> ;
  wire \adder_4bit_15.a<2> ;
  wire \adder_4bit_15.a<3> ;
  wire \adder_4bit_15.b<0> ;
  wire \adder_4bit_15.b<1> ;
  wire \adder_4bit_15.b<2> ;
  wire \adder_4bit_15.b<3> ;
  wire \adder_4bit_15.c<0> ;
  wire \adder_4bit_15.c<1> ;
  wire \adder_4bit_15.c<2> ;
  wire \adder_4bit_15.c<3> ;
  wire \adder_4bit_15.s<0> ;
  wire \adder_4bit_15.s<1> ;
  wire \adder_4bit_15.s<2> ;
  wire \adder_4bit_15.s<3> ;
  wire \adder_4bit_15.s<4> ;
  wire \adder_4bit_15.sign ;
  wire \adder_4bit_16.a<0> ;
  wire \adder_4bit_16.a<1> ;
  wire \adder_4bit_16.a<2> ;
  wire \adder_4bit_16.a<3> ;
  wire \adder_4bit_16.b<0> ;
  wire \adder_4bit_16.b<1> ;
  wire \adder_4bit_16.b<2> ;
  wire \adder_4bit_16.b<3> ;
  wire \adder_4bit_16.c<0> ;
  wire \adder_4bit_16.c<1> ;
  wire \adder_4bit_16.c<2> ;
  wire \adder_4bit_16.c<3> ;
  wire \adder_4bit_16.s<0> ;
  wire \adder_4bit_16.s<1> ;
  wire \adder_4bit_16.s<2> ;
  wire \adder_4bit_16.s<3> ;
  wire \adder_4bit_16.s<4> ;
  wire \adder_4bit_16.sign ;
  wire \adder_4bit_17.a<0> ;
  wire \adder_4bit_17.a<1> ;
  wire \adder_4bit_17.a<2> ;
  wire \adder_4bit_17.a<3> ;
  wire \adder_4bit_17.b<0> ;
  wire \adder_4bit_17.b<1> ;
  wire \adder_4bit_17.b<2> ;
  wire \adder_4bit_17.b<3> ;
  wire \adder_4bit_17.c<0> ;
  wire \adder_4bit_17.c<1> ;
  wire \adder_4bit_17.c<2> ;
  wire \adder_4bit_17.c<3> ;
  wire \adder_4bit_17.s<0> ;
  wire \adder_4bit_17.s<1> ;
  wire \adder_4bit_17.s<2> ;
  wire \adder_4bit_17.s<3> ;
  wire \adder_4bit_17.s<4> ;
  wire \adder_4bit_17.sign ;
  wire \adder_4bit_18.a<0> ;
  wire \adder_4bit_18.a<1> ;
  wire \adder_4bit_18.a<2> ;
  wire \adder_4bit_18.a<3> ;
  wire \adder_4bit_18.b<0> ;
  wire \adder_4bit_18.b<1> ;
  wire \adder_4bit_18.b<2> ;
  wire \adder_4bit_18.b<3> ;
  wire \adder_4bit_18.c<0> ;
  wire \adder_4bit_18.c<1> ;
  wire \adder_4bit_18.c<2> ;
  wire \adder_4bit_18.c<3> ;
  wire \adder_4bit_18.s<0> ;
  wire \adder_4bit_18.s<1> ;
  wire \adder_4bit_18.s<2> ;
  wire \adder_4bit_18.s<3> ;
  wire \adder_4bit_18.s<4> ;
  wire \adder_4bit_18.sign ;
  wire \adder_4bit_19.a<0> ;
  wire \adder_4bit_19.a<1> ;
  wire \adder_4bit_19.a<2> ;
  wire \adder_4bit_19.a<3> ;
  wire \adder_4bit_19.b<0> ;
  wire \adder_4bit_19.b<1> ;
  wire \adder_4bit_19.b<2> ;
  wire \adder_4bit_19.b<3> ;
  wire \adder_4bit_19.c<0> ;
  wire \adder_4bit_19.c<1> ;
  wire \adder_4bit_19.c<2> ;
  wire \adder_4bit_19.c<3> ;
  wire \adder_4bit_19.s<0> ;
  wire \adder_4bit_19.s<1> ;
  wire \adder_4bit_19.s<2> ;
  wire \adder_4bit_19.s<3> ;
  wire \adder_4bit_19.s<4> ;
  wire \adder_4bit_19.sign ;
  wire \adder_4bit_2.a<0> ;
  wire \adder_4bit_2.a<1> ;
  wire \adder_4bit_2.a<2> ;
  wire \adder_4bit_2.a<3> ;
  wire \adder_4bit_2.b<0> ;
  wire \adder_4bit_2.b<1> ;
  wire \adder_4bit_2.b<2> ;
  wire \adder_4bit_2.b<3> ;
  wire \adder_4bit_2.c<0> ;
  wire \adder_4bit_2.c<1> ;
  wire \adder_4bit_2.c<2> ;
  wire \adder_4bit_2.c<3> ;
  wire \adder_4bit_2.s<0> ;
  wire \adder_4bit_2.s<1> ;
  wire \adder_4bit_2.s<2> ;
  wire \adder_4bit_2.s<3> ;
  wire \adder_4bit_2.s<4> ;
  wire \adder_4bit_2.sign ;
  wire \adder_4bit_20.a<0> ;
  wire \adder_4bit_20.a<1> ;
  wire \adder_4bit_20.a<2> ;
  wire \adder_4bit_20.a<3> ;
  wire \adder_4bit_20.b<0> ;
  wire \adder_4bit_20.b<1> ;
  wire \adder_4bit_20.b<2> ;
  wire \adder_4bit_20.b<3> ;
  wire \adder_4bit_20.c<0> ;
  wire \adder_4bit_20.c<1> ;
  wire \adder_4bit_20.c<2> ;
  wire \adder_4bit_20.c<3> ;
  wire \adder_4bit_20.s<0> ;
  wire \adder_4bit_20.s<1> ;
  wire \adder_4bit_20.s<2> ;
  wire \adder_4bit_20.s<3> ;
  wire \adder_4bit_20.s<4> ;
  wire \adder_4bit_20.sign ;
  wire \adder_4bit_21.a<0> ;
  wire \adder_4bit_21.a<1> ;
  wire \adder_4bit_21.a<2> ;
  wire \adder_4bit_21.a<3> ;
  wire \adder_4bit_21.b<0> ;
  wire \adder_4bit_21.b<1> ;
  wire \adder_4bit_21.b<2> ;
  wire \adder_4bit_21.b<3> ;
  wire \adder_4bit_21.c<0> ;
  wire \adder_4bit_21.c<1> ;
  wire \adder_4bit_21.c<2> ;
  wire \adder_4bit_21.c<3> ;
  wire \adder_4bit_21.s<0> ;
  wire \adder_4bit_21.s<1> ;
  wire \adder_4bit_21.s<2> ;
  wire \adder_4bit_21.s<3> ;
  wire \adder_4bit_21.s<4> ;
  wire \adder_4bit_21.sign ;
  wire \adder_4bit_22.a<0> ;
  wire \adder_4bit_22.a<1> ;
  wire \adder_4bit_22.a<2> ;
  wire \adder_4bit_22.a<3> ;
  wire \adder_4bit_22.b<0> ;
  wire \adder_4bit_22.b<1> ;
  wire \adder_4bit_22.b<2> ;
  wire \adder_4bit_22.b<3> ;
  wire \adder_4bit_22.c<0> ;
  wire \adder_4bit_22.c<1> ;
  wire \adder_4bit_22.c<2> ;
  wire \adder_4bit_22.c<3> ;
  wire \adder_4bit_22.s<0> ;
  wire \adder_4bit_22.s<1> ;
  wire \adder_4bit_22.s<2> ;
  wire \adder_4bit_22.s<3> ;
  wire \adder_4bit_22.s<4> ;
  wire \adder_4bit_22.sign ;
  wire \adder_4bit_23.a<0> ;
  wire \adder_4bit_23.a<1> ;
  wire \adder_4bit_23.a<2> ;
  wire \adder_4bit_23.a<3> ;
  wire \adder_4bit_23.b<0> ;
  wire \adder_4bit_23.b<1> ;
  wire \adder_4bit_23.b<2> ;
  wire \adder_4bit_23.b<3> ;
  wire \adder_4bit_23.c<0> ;
  wire \adder_4bit_23.c<1> ;
  wire \adder_4bit_23.c<2> ;
  wire \adder_4bit_23.c<3> ;
  wire \adder_4bit_23.s<0> ;
  wire \adder_4bit_23.s<1> ;
  wire \adder_4bit_23.s<2> ;
  wire \adder_4bit_23.s<3> ;
  wire \adder_4bit_23.s<4> ;
  wire \adder_4bit_23.sign ;
  wire \adder_4bit_24.a<0> ;
  wire \adder_4bit_24.a<1> ;
  wire \adder_4bit_24.a<2> ;
  wire \adder_4bit_24.a<3> ;
  wire \adder_4bit_24.b<0> ;
  wire \adder_4bit_24.b<1> ;
  wire \adder_4bit_24.b<2> ;
  wire \adder_4bit_24.b<3> ;
  wire \adder_4bit_24.c<0> ;
  wire \adder_4bit_24.c<1> ;
  wire \adder_4bit_24.c<2> ;
  wire \adder_4bit_24.c<3> ;
  wire \adder_4bit_24.s<0> ;
  wire \adder_4bit_24.s<1> ;
  wire \adder_4bit_24.s<2> ;
  wire \adder_4bit_24.s<3> ;
  wire \adder_4bit_24.s<4> ;
  wire \adder_4bit_24.sign ;
  wire \adder_4bit_25.a<0> ;
  wire \adder_4bit_25.a<1> ;
  wire \adder_4bit_25.a<2> ;
  wire \adder_4bit_25.a<3> ;
  wire \adder_4bit_25.b<0> ;
  wire \adder_4bit_25.b<1> ;
  wire \adder_4bit_25.b<2> ;
  wire \adder_4bit_25.b<3> ;
  wire \adder_4bit_25.c<0> ;
  wire \adder_4bit_25.c<1> ;
  wire \adder_4bit_25.c<2> ;
  wire \adder_4bit_25.c<3> ;
  wire \adder_4bit_25.s<0> ;
  wire \adder_4bit_25.s<1> ;
  wire \adder_4bit_25.s<2> ;
  wire \adder_4bit_25.s<3> ;
  wire \adder_4bit_25.s<4> ;
  wire \adder_4bit_25.sign ;
  wire \adder_4bit_26.a<0> ;
  wire \adder_4bit_26.a<1> ;
  wire \adder_4bit_26.a<2> ;
  wire \adder_4bit_26.a<3> ;
  wire \adder_4bit_26.b<0> ;
  wire \adder_4bit_26.b<1> ;
  wire \adder_4bit_26.b<2> ;
  wire \adder_4bit_26.b<3> ;
  wire \adder_4bit_26.c<0> ;
  wire \adder_4bit_26.c<1> ;
  wire \adder_4bit_26.c<2> ;
  wire \adder_4bit_26.c<3> ;
  wire \adder_4bit_26.s<0> ;
  wire \adder_4bit_26.s<1> ;
  wire \adder_4bit_26.s<2> ;
  wire \adder_4bit_26.s<3> ;
  wire \adder_4bit_26.s<4> ;
  wire \adder_4bit_26.sign ;
  wire \adder_4bit_27.a<0> ;
  wire \adder_4bit_27.a<1> ;
  wire \adder_4bit_27.a<2> ;
  wire \adder_4bit_27.a<3> ;
  wire \adder_4bit_27.b<0> ;
  wire \adder_4bit_27.b<1> ;
  wire \adder_4bit_27.b<2> ;
  wire \adder_4bit_27.b<3> ;
  wire \adder_4bit_27.c<0> ;
  wire \adder_4bit_27.c<1> ;
  wire \adder_4bit_27.c<2> ;
  wire \adder_4bit_27.c<3> ;
  wire \adder_4bit_27.s<0> ;
  wire \adder_4bit_27.s<1> ;
  wire \adder_4bit_27.s<2> ;
  wire \adder_4bit_27.s<3> ;
  wire \adder_4bit_27.s<4> ;
  wire \adder_4bit_27.sign ;
  wire \adder_4bit_28.a<0> ;
  wire \adder_4bit_28.a<1> ;
  wire \adder_4bit_28.a<2> ;
  wire \adder_4bit_28.a<3> ;
  wire \adder_4bit_28.b<0> ;
  wire \adder_4bit_28.b<1> ;
  wire \adder_4bit_28.b<2> ;
  wire \adder_4bit_28.b<3> ;
  wire \adder_4bit_28.c<0> ;
  wire \adder_4bit_28.c<1> ;
  wire \adder_4bit_28.c<2> ;
  wire \adder_4bit_28.c<3> ;
  wire \adder_4bit_28.s<0> ;
  wire \adder_4bit_28.s<1> ;
  wire \adder_4bit_28.s<2> ;
  wire \adder_4bit_28.s<3> ;
  wire \adder_4bit_28.s<4> ;
  wire \adder_4bit_28.sign ;
  wire \adder_4bit_29.a<0> ;
  wire \adder_4bit_29.a<1> ;
  wire \adder_4bit_29.a<2> ;
  wire \adder_4bit_29.a<3> ;
  wire \adder_4bit_29.b<0> ;
  wire \adder_4bit_29.b<1> ;
  wire \adder_4bit_29.b<2> ;
  wire \adder_4bit_29.b<3> ;
  wire \adder_4bit_29.c<0> ;
  wire \adder_4bit_29.c<1> ;
  wire \adder_4bit_29.c<2> ;
  wire \adder_4bit_29.c<3> ;
  wire \adder_4bit_29.s<0> ;
  wire \adder_4bit_29.s<1> ;
  wire \adder_4bit_29.s<2> ;
  wire \adder_4bit_29.s<3> ;
  wire \adder_4bit_29.s<4> ;
  wire \adder_4bit_29.sign ;
  wire \adder_4bit_3.a<0> ;
  wire \adder_4bit_3.a<1> ;
  wire \adder_4bit_3.a<2> ;
  wire \adder_4bit_3.a<3> ;
  wire \adder_4bit_3.b<0> ;
  wire \adder_4bit_3.b<1> ;
  wire \adder_4bit_3.b<2> ;
  wire \adder_4bit_3.b<3> ;
  wire \adder_4bit_3.c<0> ;
  wire \adder_4bit_3.c<1> ;
  wire \adder_4bit_3.c<2> ;
  wire \adder_4bit_3.c<3> ;
  wire \adder_4bit_3.s<0> ;
  wire \adder_4bit_3.s<1> ;
  wire \adder_4bit_3.s<2> ;
  wire \adder_4bit_3.s<3> ;
  wire \adder_4bit_3.s<4> ;
  wire \adder_4bit_3.sign ;
  wire \adder_4bit_30.a<0> ;
  wire \adder_4bit_30.a<1> ;
  wire \adder_4bit_30.a<2> ;
  wire \adder_4bit_30.a<3> ;
  wire \adder_4bit_30.b<0> ;
  wire \adder_4bit_30.b<1> ;
  wire \adder_4bit_30.b<2> ;
  wire \adder_4bit_30.b<3> ;
  wire \adder_4bit_30.c<0> ;
  wire \adder_4bit_30.c<1> ;
  wire \adder_4bit_30.c<2> ;
  wire \adder_4bit_30.c<3> ;
  wire \adder_4bit_30.s<0> ;
  wire \adder_4bit_30.s<1> ;
  wire \adder_4bit_30.s<2> ;
  wire \adder_4bit_30.s<3> ;
  wire \adder_4bit_30.s<4> ;
  wire \adder_4bit_30.sign ;
  wire \adder_4bit_31.a<0> ;
  wire \adder_4bit_31.a<1> ;
  wire \adder_4bit_31.a<2> ;
  wire \adder_4bit_31.a<3> ;
  wire \adder_4bit_31.b<0> ;
  wire \adder_4bit_31.b<1> ;
  wire \adder_4bit_31.b<2> ;
  wire \adder_4bit_31.b<3> ;
  wire \adder_4bit_31.c<0> ;
  wire \adder_4bit_31.c<1> ;
  wire \adder_4bit_31.c<2> ;
  wire \adder_4bit_31.c<3> ;
  wire \adder_4bit_31.s<0> ;
  wire \adder_4bit_31.s<1> ;
  wire \adder_4bit_31.s<2> ;
  wire \adder_4bit_31.s<3> ;
  wire \adder_4bit_31.s<4> ;
  wire \adder_4bit_31.sign ;
  wire \adder_4bit_4.a<0> ;
  wire \adder_4bit_4.a<1> ;
  wire \adder_4bit_4.a<2> ;
  wire \adder_4bit_4.a<3> ;
  wire \adder_4bit_4.b<0> ;
  wire \adder_4bit_4.b<1> ;
  wire \adder_4bit_4.b<2> ;
  wire \adder_4bit_4.b<3> ;
  wire \adder_4bit_4.c<0> ;
  wire \adder_4bit_4.c<1> ;
  wire \adder_4bit_4.c<2> ;
  wire \adder_4bit_4.c<3> ;
  wire \adder_4bit_4.s<0> ;
  wire \adder_4bit_4.s<1> ;
  wire \adder_4bit_4.s<2> ;
  wire \adder_4bit_4.s<3> ;
  wire \adder_4bit_4.s<4> ;
  wire \adder_4bit_4.sign ;
  wire \adder_4bit_5.a<0> ;
  wire \adder_4bit_5.a<1> ;
  wire \adder_4bit_5.a<2> ;
  wire \adder_4bit_5.a<3> ;
  wire \adder_4bit_5.b<0> ;
  wire \adder_4bit_5.b<1> ;
  wire \adder_4bit_5.b<2> ;
  wire \adder_4bit_5.b<3> ;
  wire \adder_4bit_5.c<0> ;
  wire \adder_4bit_5.c<1> ;
  wire \adder_4bit_5.c<2> ;
  wire \adder_4bit_5.c<3> ;
  wire \adder_4bit_5.s<0> ;
  wire \adder_4bit_5.s<1> ;
  wire \adder_4bit_5.s<2> ;
  wire \adder_4bit_5.s<3> ;
  wire \adder_4bit_5.s<4> ;
  wire \adder_4bit_5.sign ;
  wire \adder_4bit_6.a<0> ;
  wire \adder_4bit_6.a<1> ;
  wire \adder_4bit_6.a<2> ;
  wire \adder_4bit_6.a<3> ;
  wire \adder_4bit_6.b<0> ;
  wire \adder_4bit_6.b<1> ;
  wire \adder_4bit_6.b<2> ;
  wire \adder_4bit_6.b<3> ;
  wire \adder_4bit_6.c<0> ;
  wire \adder_4bit_6.c<1> ;
  wire \adder_4bit_6.c<2> ;
  wire \adder_4bit_6.c<3> ;
  wire \adder_4bit_6.s<0> ;
  wire \adder_4bit_6.s<1> ;
  wire \adder_4bit_6.s<2> ;
  wire \adder_4bit_6.s<3> ;
  wire \adder_4bit_6.s<4> ;
  wire \adder_4bit_6.sign ;
  wire \adder_4bit_7.a<0> ;
  wire \adder_4bit_7.a<1> ;
  wire \adder_4bit_7.a<2> ;
  wire \adder_4bit_7.a<3> ;
  wire \adder_4bit_7.b<0> ;
  wire \adder_4bit_7.b<1> ;
  wire \adder_4bit_7.b<2> ;
  wire \adder_4bit_7.b<3> ;
  wire \adder_4bit_7.c<0> ;
  wire \adder_4bit_7.c<1> ;
  wire \adder_4bit_7.c<2> ;
  wire \adder_4bit_7.c<3> ;
  wire \adder_4bit_7.s<0> ;
  wire \adder_4bit_7.s<1> ;
  wire \adder_4bit_7.s<2> ;
  wire \adder_4bit_7.s<3> ;
  wire \adder_4bit_7.s<4> ;
  wire \adder_4bit_7.sign ;
  wire \adder_4bit_8.a<0> ;
  wire \adder_4bit_8.a<1> ;
  wire \adder_4bit_8.a<2> ;
  wire \adder_4bit_8.a<3> ;
  wire \adder_4bit_8.b<0> ;
  wire \adder_4bit_8.b<1> ;
  wire \adder_4bit_8.b<2> ;
  wire \adder_4bit_8.b<3> ;
  wire \adder_4bit_8.c<0> ;
  wire \adder_4bit_8.c<1> ;
  wire \adder_4bit_8.c<2> ;
  wire \adder_4bit_8.c<3> ;
  wire \adder_4bit_8.s<0> ;
  wire \adder_4bit_8.s<1> ;
  wire \adder_4bit_8.s<2> ;
  wire \adder_4bit_8.s<3> ;
  wire \adder_4bit_8.s<4> ;
  wire \adder_4bit_8.sign ;
  wire \adder_4bit_9.a<0> ;
  wire \adder_4bit_9.a<1> ;
  wire \adder_4bit_9.a<2> ;
  wire \adder_4bit_9.a<3> ;
  wire \adder_4bit_9.b<0> ;
  wire \adder_4bit_9.b<1> ;
  wire \adder_4bit_9.b<2> ;
  wire \adder_4bit_9.b<3> ;
  wire \adder_4bit_9.c<0> ;
  wire \adder_4bit_9.c<1> ;
  wire \adder_4bit_9.c<2> ;
  wire \adder_4bit_9.c<3> ;
  wire \adder_4bit_9.s<0> ;
  wire \adder_4bit_9.s<1> ;
  wire \adder_4bit_9.s<2> ;
  wire \adder_4bit_9.s<3> ;
  wire \adder_4bit_9.s<4> ;
  wire \adder_4bit_9.sign ;
  wire \adder_5bit_0.a<0> ;
  wire \adder_5bit_0.a<1> ;
  wire \adder_5bit_0.a<2> ;
  wire \adder_5bit_0.a<3> ;
  wire \adder_5bit_0.a<4> ;
  wire \adder_5bit_0.b<0> ;
  wire \adder_5bit_0.b<1> ;
  wire \adder_5bit_0.b<2> ;
  wire \adder_5bit_0.b<3> ;
  wire \adder_5bit_0.b<4> ;
  wire \adder_5bit_0.c<0> ;
  wire \adder_5bit_0.c<1> ;
  wire \adder_5bit_0.c<2> ;
  wire \adder_5bit_0.c<3> ;
  wire \adder_5bit_0.c<4> ;
  wire \adder_5bit_0.s<0> ;
  wire \adder_5bit_0.s<1> ;
  wire \adder_5bit_0.s<2> ;
  wire \adder_5bit_0.s<3> ;
  wire \adder_5bit_0.s<4> ;
  wire \adder_5bit_0.s<5> ;
  wire \adder_5bit_0.sign ;
  wire \adder_5bit_1.a<0> ;
  wire \adder_5bit_1.a<1> ;
  wire \adder_5bit_1.a<2> ;
  wire \adder_5bit_1.a<3> ;
  wire \adder_5bit_1.a<4> ;
  wire \adder_5bit_1.b<0> ;
  wire \adder_5bit_1.b<1> ;
  wire \adder_5bit_1.b<2> ;
  wire \adder_5bit_1.b<3> ;
  wire \adder_5bit_1.b<4> ;
  wire \adder_5bit_1.c<0> ;
  wire \adder_5bit_1.c<1> ;
  wire \adder_5bit_1.c<2> ;
  wire \adder_5bit_1.c<3> ;
  wire \adder_5bit_1.c<4> ;
  wire \adder_5bit_1.s<0> ;
  wire \adder_5bit_1.s<1> ;
  wire \adder_5bit_1.s<2> ;
  wire \adder_5bit_1.s<3> ;
  wire \adder_5bit_1.s<4> ;
  wire \adder_5bit_1.s<5> ;
  wire \adder_5bit_1.sign ;
  wire \adder_5bit_10.a<0> ;
  wire \adder_5bit_10.a<1> ;
  wire \adder_5bit_10.a<2> ;
  wire \adder_5bit_10.a<3> ;
  wire \adder_5bit_10.a<4> ;
  wire \adder_5bit_10.b<0> ;
  wire \adder_5bit_10.b<1> ;
  wire \adder_5bit_10.b<2> ;
  wire \adder_5bit_10.b<3> ;
  wire \adder_5bit_10.b<4> ;
  wire \adder_5bit_10.c<0> ;
  wire \adder_5bit_10.c<1> ;
  wire \adder_5bit_10.c<2> ;
  wire \adder_5bit_10.c<3> ;
  wire \adder_5bit_10.c<4> ;
  wire \adder_5bit_10.s<0> ;
  wire \adder_5bit_10.s<1> ;
  wire \adder_5bit_10.s<2> ;
  wire \adder_5bit_10.s<3> ;
  wire \adder_5bit_10.s<4> ;
  wire \adder_5bit_10.s<5> ;
  wire \adder_5bit_10.sign ;
  wire \adder_5bit_11.a<0> ;
  wire \adder_5bit_11.a<1> ;
  wire \adder_5bit_11.a<2> ;
  wire \adder_5bit_11.a<3> ;
  wire \adder_5bit_11.a<4> ;
  wire \adder_5bit_11.b<0> ;
  wire \adder_5bit_11.b<1> ;
  wire \adder_5bit_11.b<2> ;
  wire \adder_5bit_11.b<3> ;
  wire \adder_5bit_11.b<4> ;
  wire \adder_5bit_11.c<0> ;
  wire \adder_5bit_11.c<1> ;
  wire \adder_5bit_11.c<2> ;
  wire \adder_5bit_11.c<3> ;
  wire \adder_5bit_11.c<4> ;
  wire \adder_5bit_11.s<0> ;
  wire \adder_5bit_11.s<1> ;
  wire \adder_5bit_11.s<2> ;
  wire \adder_5bit_11.s<3> ;
  wire \adder_5bit_11.s<4> ;
  wire \adder_5bit_11.s<5> ;
  wire \adder_5bit_11.sign ;
  wire \adder_5bit_12.a<0> ;
  wire \adder_5bit_12.a<1> ;
  wire \adder_5bit_12.a<2> ;
  wire \adder_5bit_12.a<3> ;
  wire \adder_5bit_12.a<4> ;
  wire \adder_5bit_12.b<0> ;
  wire \adder_5bit_12.b<1> ;
  wire \adder_5bit_12.b<2> ;
  wire \adder_5bit_12.b<3> ;
  wire \adder_5bit_12.b<4> ;
  wire \adder_5bit_12.c<0> ;
  wire \adder_5bit_12.c<1> ;
  wire \adder_5bit_12.c<2> ;
  wire \adder_5bit_12.c<3> ;
  wire \adder_5bit_12.c<4> ;
  wire \adder_5bit_12.s<0> ;
  wire \adder_5bit_12.s<1> ;
  wire \adder_5bit_12.s<2> ;
  wire \adder_5bit_12.s<3> ;
  wire \adder_5bit_12.s<4> ;
  wire \adder_5bit_12.s<5> ;
  wire \adder_5bit_12.sign ;
  wire \adder_5bit_13.a<0> ;
  wire \adder_5bit_13.a<1> ;
  wire \adder_5bit_13.a<2> ;
  wire \adder_5bit_13.a<3> ;
  wire \adder_5bit_13.a<4> ;
  wire \adder_5bit_13.b<0> ;
  wire \adder_5bit_13.b<1> ;
  wire \adder_5bit_13.b<2> ;
  wire \adder_5bit_13.b<3> ;
  wire \adder_5bit_13.b<4> ;
  wire \adder_5bit_13.c<0> ;
  wire \adder_5bit_13.c<1> ;
  wire \adder_5bit_13.c<2> ;
  wire \adder_5bit_13.c<3> ;
  wire \adder_5bit_13.c<4> ;
  wire \adder_5bit_13.s<0> ;
  wire \adder_5bit_13.s<1> ;
  wire \adder_5bit_13.s<2> ;
  wire \adder_5bit_13.s<3> ;
  wire \adder_5bit_13.s<4> ;
  wire \adder_5bit_13.s<5> ;
  wire \adder_5bit_13.sign ;
  wire \adder_5bit_14.a<0> ;
  wire \adder_5bit_14.a<1> ;
  wire \adder_5bit_14.a<2> ;
  wire \adder_5bit_14.a<3> ;
  wire \adder_5bit_14.a<4> ;
  wire \adder_5bit_14.b<0> ;
  wire \adder_5bit_14.b<1> ;
  wire \adder_5bit_14.b<2> ;
  wire \adder_5bit_14.b<3> ;
  wire \adder_5bit_14.b<4> ;
  wire \adder_5bit_14.c<0> ;
  wire \adder_5bit_14.c<1> ;
  wire \adder_5bit_14.c<2> ;
  wire \adder_5bit_14.c<3> ;
  wire \adder_5bit_14.c<4> ;
  wire \adder_5bit_14.s<0> ;
  wire \adder_5bit_14.s<1> ;
  wire \adder_5bit_14.s<2> ;
  wire \adder_5bit_14.s<3> ;
  wire \adder_5bit_14.s<4> ;
  wire \adder_5bit_14.s<5> ;
  wire \adder_5bit_14.sign ;
  wire \adder_5bit_15.a<0> ;
  wire \adder_5bit_15.a<1> ;
  wire \adder_5bit_15.a<2> ;
  wire \adder_5bit_15.a<3> ;
  wire \adder_5bit_15.a<4> ;
  wire \adder_5bit_15.b<0> ;
  wire \adder_5bit_15.b<1> ;
  wire \adder_5bit_15.b<2> ;
  wire \adder_5bit_15.b<3> ;
  wire \adder_5bit_15.b<4> ;
  wire \adder_5bit_15.c<0> ;
  wire \adder_5bit_15.c<1> ;
  wire \adder_5bit_15.c<2> ;
  wire \adder_5bit_15.c<3> ;
  wire \adder_5bit_15.c<4> ;
  wire \adder_5bit_15.s<0> ;
  wire \adder_5bit_15.s<1> ;
  wire \adder_5bit_15.s<2> ;
  wire \adder_5bit_15.s<3> ;
  wire \adder_5bit_15.s<4> ;
  wire \adder_5bit_15.s<5> ;
  wire \adder_5bit_15.sign ;
  wire \adder_5bit_2.a<0> ;
  wire \adder_5bit_2.a<1> ;
  wire \adder_5bit_2.a<2> ;
  wire \adder_5bit_2.a<3> ;
  wire \adder_5bit_2.a<4> ;
  wire \adder_5bit_2.b<0> ;
  wire \adder_5bit_2.b<1> ;
  wire \adder_5bit_2.b<2> ;
  wire \adder_5bit_2.b<3> ;
  wire \adder_5bit_2.b<4> ;
  wire \adder_5bit_2.c<0> ;
  wire \adder_5bit_2.c<1> ;
  wire \adder_5bit_2.c<2> ;
  wire \adder_5bit_2.c<3> ;
  wire \adder_5bit_2.c<4> ;
  wire \adder_5bit_2.s<0> ;
  wire \adder_5bit_2.s<1> ;
  wire \adder_5bit_2.s<2> ;
  wire \adder_5bit_2.s<3> ;
  wire \adder_5bit_2.s<4> ;
  wire \adder_5bit_2.s<5> ;
  wire \adder_5bit_2.sign ;
  wire \adder_5bit_3.a<0> ;
  wire \adder_5bit_3.a<1> ;
  wire \adder_5bit_3.a<2> ;
  wire \adder_5bit_3.a<3> ;
  wire \adder_5bit_3.a<4> ;
  wire \adder_5bit_3.b<0> ;
  wire \adder_5bit_3.b<1> ;
  wire \adder_5bit_3.b<2> ;
  wire \adder_5bit_3.b<3> ;
  wire \adder_5bit_3.b<4> ;
  wire \adder_5bit_3.c<0> ;
  wire \adder_5bit_3.c<1> ;
  wire \adder_5bit_3.c<2> ;
  wire \adder_5bit_3.c<3> ;
  wire \adder_5bit_3.c<4> ;
  wire \adder_5bit_3.s<0> ;
  wire \adder_5bit_3.s<1> ;
  wire \adder_5bit_3.s<2> ;
  wire \adder_5bit_3.s<3> ;
  wire \adder_5bit_3.s<4> ;
  wire \adder_5bit_3.s<5> ;
  wire \adder_5bit_3.sign ;
  wire \adder_5bit_4.a<0> ;
  wire \adder_5bit_4.a<1> ;
  wire \adder_5bit_4.a<2> ;
  wire \adder_5bit_4.a<3> ;
  wire \adder_5bit_4.a<4> ;
  wire \adder_5bit_4.b<0> ;
  wire \adder_5bit_4.b<1> ;
  wire \adder_5bit_4.b<2> ;
  wire \adder_5bit_4.b<3> ;
  wire \adder_5bit_4.b<4> ;
  wire \adder_5bit_4.c<0> ;
  wire \adder_5bit_4.c<1> ;
  wire \adder_5bit_4.c<2> ;
  wire \adder_5bit_4.c<3> ;
  wire \adder_5bit_4.c<4> ;
  wire \adder_5bit_4.s<0> ;
  wire \adder_5bit_4.s<1> ;
  wire \adder_5bit_4.s<2> ;
  wire \adder_5bit_4.s<3> ;
  wire \adder_5bit_4.s<4> ;
  wire \adder_5bit_4.s<5> ;
  wire \adder_5bit_4.sign ;
  wire \adder_5bit_5.a<0> ;
  wire \adder_5bit_5.a<1> ;
  wire \adder_5bit_5.a<2> ;
  wire \adder_5bit_5.a<3> ;
  wire \adder_5bit_5.a<4> ;
  wire \adder_5bit_5.b<0> ;
  wire \adder_5bit_5.b<1> ;
  wire \adder_5bit_5.b<2> ;
  wire \adder_5bit_5.b<3> ;
  wire \adder_5bit_5.b<4> ;
  wire \adder_5bit_5.c<0> ;
  wire \adder_5bit_5.c<1> ;
  wire \adder_5bit_5.c<2> ;
  wire \adder_5bit_5.c<3> ;
  wire \adder_5bit_5.c<4> ;
  wire \adder_5bit_5.s<0> ;
  wire \adder_5bit_5.s<1> ;
  wire \adder_5bit_5.s<2> ;
  wire \adder_5bit_5.s<3> ;
  wire \adder_5bit_5.s<4> ;
  wire \adder_5bit_5.s<5> ;
  wire \adder_5bit_5.sign ;
  wire \adder_5bit_6.a<0> ;
  wire \adder_5bit_6.a<1> ;
  wire \adder_5bit_6.a<2> ;
  wire \adder_5bit_6.a<3> ;
  wire \adder_5bit_6.a<4> ;
  wire \adder_5bit_6.b<0> ;
  wire \adder_5bit_6.b<1> ;
  wire \adder_5bit_6.b<2> ;
  wire \adder_5bit_6.b<3> ;
  wire \adder_5bit_6.b<4> ;
  wire \adder_5bit_6.c<0> ;
  wire \adder_5bit_6.c<1> ;
  wire \adder_5bit_6.c<2> ;
  wire \adder_5bit_6.c<3> ;
  wire \adder_5bit_6.c<4> ;
  wire \adder_5bit_6.s<0> ;
  wire \adder_5bit_6.s<1> ;
  wire \adder_5bit_6.s<2> ;
  wire \adder_5bit_6.s<3> ;
  wire \adder_5bit_6.s<4> ;
  wire \adder_5bit_6.s<5> ;
  wire \adder_5bit_6.sign ;
  wire \adder_5bit_7.a<0> ;
  wire \adder_5bit_7.a<1> ;
  wire \adder_5bit_7.a<2> ;
  wire \adder_5bit_7.a<3> ;
  wire \adder_5bit_7.a<4> ;
  wire \adder_5bit_7.b<0> ;
  wire \adder_5bit_7.b<1> ;
  wire \adder_5bit_7.b<2> ;
  wire \adder_5bit_7.b<3> ;
  wire \adder_5bit_7.b<4> ;
  wire \adder_5bit_7.c<0> ;
  wire \adder_5bit_7.c<1> ;
  wire \adder_5bit_7.c<2> ;
  wire \adder_5bit_7.c<3> ;
  wire \adder_5bit_7.c<4> ;
  wire \adder_5bit_7.s<0> ;
  wire \adder_5bit_7.s<1> ;
  wire \adder_5bit_7.s<2> ;
  wire \adder_5bit_7.s<3> ;
  wire \adder_5bit_7.s<4> ;
  wire \adder_5bit_7.s<5> ;
  wire \adder_5bit_7.sign ;
  wire \adder_5bit_8.a<0> ;
  wire \adder_5bit_8.a<1> ;
  wire \adder_5bit_8.a<2> ;
  wire \adder_5bit_8.a<3> ;
  wire \adder_5bit_8.a<4> ;
  wire \adder_5bit_8.b<0> ;
  wire \adder_5bit_8.b<1> ;
  wire \adder_5bit_8.b<2> ;
  wire \adder_5bit_8.b<3> ;
  wire \adder_5bit_8.b<4> ;
  wire \adder_5bit_8.c<0> ;
  wire \adder_5bit_8.c<1> ;
  wire \adder_5bit_8.c<2> ;
  wire \adder_5bit_8.c<3> ;
  wire \adder_5bit_8.c<4> ;
  wire \adder_5bit_8.s<0> ;
  wire \adder_5bit_8.s<1> ;
  wire \adder_5bit_8.s<2> ;
  wire \adder_5bit_8.s<3> ;
  wire \adder_5bit_8.s<4> ;
  wire \adder_5bit_8.s<5> ;
  wire \adder_5bit_8.sign ;
  wire \adder_5bit_9.a<0> ;
  wire \adder_5bit_9.a<1> ;
  wire \adder_5bit_9.a<2> ;
  wire \adder_5bit_9.a<3> ;
  wire \adder_5bit_9.a<4> ;
  wire \adder_5bit_9.b<0> ;
  wire \adder_5bit_9.b<1> ;
  wire \adder_5bit_9.b<2> ;
  wire \adder_5bit_9.b<3> ;
  wire \adder_5bit_9.b<4> ;
  wire \adder_5bit_9.c<0> ;
  wire \adder_5bit_9.c<1> ;
  wire \adder_5bit_9.c<2> ;
  wire \adder_5bit_9.c<3> ;
  wire \adder_5bit_9.c<4> ;
  wire \adder_5bit_9.s<0> ;
  wire \adder_5bit_9.s<1> ;
  wire \adder_5bit_9.s<2> ;
  wire \adder_5bit_9.s<3> ;
  wire \adder_5bit_9.s<4> ;
  wire \adder_5bit_9.s<5> ;
  wire \adder_5bit_9.sign ;
  wire \adder_6bit_0.a<0> ;
  wire \adder_6bit_0.a<1> ;
  wire \adder_6bit_0.a<2> ;
  wire \adder_6bit_0.a<3> ;
  wire \adder_6bit_0.a<4> ;
  wire \adder_6bit_0.a<5> ;
  wire \adder_6bit_0.b<0> ;
  wire \adder_6bit_0.b<1> ;
  wire \adder_6bit_0.b<2> ;
  wire \adder_6bit_0.b<3> ;
  wire \adder_6bit_0.b<4> ;
  wire \adder_6bit_0.b<5> ;
  wire \adder_6bit_0.c<0> ;
  wire \adder_6bit_0.c<1> ;
  wire \adder_6bit_0.c<2> ;
  wire \adder_6bit_0.c<3> ;
  wire \adder_6bit_0.c<4> ;
  wire \adder_6bit_0.c<5> ;
  wire \adder_6bit_0.s<0> ;
  wire \adder_6bit_0.s<1> ;
  wire \adder_6bit_0.s<2> ;
  wire \adder_6bit_0.s<3> ;
  wire \adder_6bit_0.s<4> ;
  wire \adder_6bit_0.s<5> ;
  wire \adder_6bit_0.s<6> ;
  wire \adder_6bit_0.sign ;
  wire \adder_6bit_1.a<0> ;
  wire \adder_6bit_1.a<1> ;
  wire \adder_6bit_1.a<2> ;
  wire \adder_6bit_1.a<3> ;
  wire \adder_6bit_1.a<4> ;
  wire \adder_6bit_1.a<5> ;
  wire \adder_6bit_1.b<0> ;
  wire \adder_6bit_1.b<1> ;
  wire \adder_6bit_1.b<2> ;
  wire \adder_6bit_1.b<3> ;
  wire \adder_6bit_1.b<4> ;
  wire \adder_6bit_1.b<5> ;
  wire \adder_6bit_1.c<0> ;
  wire \adder_6bit_1.c<1> ;
  wire \adder_6bit_1.c<2> ;
  wire \adder_6bit_1.c<3> ;
  wire \adder_6bit_1.c<4> ;
  wire \adder_6bit_1.c<5> ;
  wire \adder_6bit_1.s<0> ;
  wire \adder_6bit_1.s<1> ;
  wire \adder_6bit_1.s<2> ;
  wire \adder_6bit_1.s<3> ;
  wire \adder_6bit_1.s<4> ;
  wire \adder_6bit_1.s<5> ;
  wire \adder_6bit_1.s<6> ;
  wire \adder_6bit_1.sign ;
  wire \adder_6bit_2.a<0> ;
  wire \adder_6bit_2.a<1> ;
  wire \adder_6bit_2.a<2> ;
  wire \adder_6bit_2.a<3> ;
  wire \adder_6bit_2.a<4> ;
  wire \adder_6bit_2.a<5> ;
  wire \adder_6bit_2.b<0> ;
  wire \adder_6bit_2.b<1> ;
  wire \adder_6bit_2.b<2> ;
  wire \adder_6bit_2.b<3> ;
  wire \adder_6bit_2.b<4> ;
  wire \adder_6bit_2.b<5> ;
  wire \adder_6bit_2.c<0> ;
  wire \adder_6bit_2.c<1> ;
  wire \adder_6bit_2.c<2> ;
  wire \adder_6bit_2.c<3> ;
  wire \adder_6bit_2.c<4> ;
  wire \adder_6bit_2.c<5> ;
  wire \adder_6bit_2.s<0> ;
  wire \adder_6bit_2.s<1> ;
  wire \adder_6bit_2.s<2> ;
  wire \adder_6bit_2.s<3> ;
  wire \adder_6bit_2.s<4> ;
  wire \adder_6bit_2.s<5> ;
  wire \adder_6bit_2.s<6> ;
  wire \adder_6bit_2.sign ;
  wire \adder_6bit_3.a<0> ;
  wire \adder_6bit_3.a<1> ;
  wire \adder_6bit_3.a<2> ;
  wire \adder_6bit_3.a<3> ;
  wire \adder_6bit_3.a<4> ;
  wire \adder_6bit_3.a<5> ;
  wire \adder_6bit_3.b<0> ;
  wire \adder_6bit_3.b<1> ;
  wire \adder_6bit_3.b<2> ;
  wire \adder_6bit_3.b<3> ;
  wire \adder_6bit_3.b<4> ;
  wire \adder_6bit_3.b<5> ;
  wire \adder_6bit_3.c<0> ;
  wire \adder_6bit_3.c<1> ;
  wire \adder_6bit_3.c<2> ;
  wire \adder_6bit_3.c<3> ;
  wire \adder_6bit_3.c<4> ;
  wire \adder_6bit_3.c<5> ;
  wire \adder_6bit_3.s<0> ;
  wire \adder_6bit_3.s<1> ;
  wire \adder_6bit_3.s<2> ;
  wire \adder_6bit_3.s<3> ;
  wire \adder_6bit_3.s<4> ;
  wire \adder_6bit_3.s<5> ;
  wire \adder_6bit_3.s<6> ;
  wire \adder_6bit_3.sign ;
  wire \adder_6bit_4.a<0> ;
  wire \adder_6bit_4.a<1> ;
  wire \adder_6bit_4.a<2> ;
  wire \adder_6bit_4.a<3> ;
  wire \adder_6bit_4.a<4> ;
  wire \adder_6bit_4.a<5> ;
  wire \adder_6bit_4.b<0> ;
  wire \adder_6bit_4.b<1> ;
  wire \adder_6bit_4.b<2> ;
  wire \adder_6bit_4.b<3> ;
  wire \adder_6bit_4.b<4> ;
  wire \adder_6bit_4.b<5> ;
  wire \adder_6bit_4.c<0> ;
  wire \adder_6bit_4.c<1> ;
  wire \adder_6bit_4.c<2> ;
  wire \adder_6bit_4.c<3> ;
  wire \adder_6bit_4.c<4> ;
  wire \adder_6bit_4.c<5> ;
  wire \adder_6bit_4.s<0> ;
  wire \adder_6bit_4.s<1> ;
  wire \adder_6bit_4.s<2> ;
  wire \adder_6bit_4.s<3> ;
  wire \adder_6bit_4.s<4> ;
  wire \adder_6bit_4.s<5> ;
  wire \adder_6bit_4.s<6> ;
  wire \adder_6bit_4.sign ;
  wire \adder_6bit_5.a<0> ;
  wire \adder_6bit_5.a<1> ;
  wire \adder_6bit_5.a<2> ;
  wire \adder_6bit_5.a<3> ;
  wire \adder_6bit_5.a<4> ;
  wire \adder_6bit_5.a<5> ;
  wire \adder_6bit_5.b<0> ;
  wire \adder_6bit_5.b<1> ;
  wire \adder_6bit_5.b<2> ;
  wire \adder_6bit_5.b<3> ;
  wire \adder_6bit_5.b<4> ;
  wire \adder_6bit_5.b<5> ;
  wire \adder_6bit_5.c<0> ;
  wire \adder_6bit_5.c<1> ;
  wire \adder_6bit_5.c<2> ;
  wire \adder_6bit_5.c<3> ;
  wire \adder_6bit_5.c<4> ;
  wire \adder_6bit_5.c<5> ;
  wire \adder_6bit_5.s<0> ;
  wire \adder_6bit_5.s<1> ;
  wire \adder_6bit_5.s<2> ;
  wire \adder_6bit_5.s<3> ;
  wire \adder_6bit_5.s<4> ;
  wire \adder_6bit_5.s<5> ;
  wire \adder_6bit_5.s<6> ;
  wire \adder_6bit_5.sign ;
  wire \adder_6bit_6.a<0> ;
  wire \adder_6bit_6.a<1> ;
  wire \adder_6bit_6.a<2> ;
  wire \adder_6bit_6.a<3> ;
  wire \adder_6bit_6.a<4> ;
  wire \adder_6bit_6.a<5> ;
  wire \adder_6bit_6.b<0> ;
  wire \adder_6bit_6.b<1> ;
  wire \adder_6bit_6.b<2> ;
  wire \adder_6bit_6.b<3> ;
  wire \adder_6bit_6.b<4> ;
  wire \adder_6bit_6.b<5> ;
  wire \adder_6bit_6.c<0> ;
  wire \adder_6bit_6.c<1> ;
  wire \adder_6bit_6.c<2> ;
  wire \adder_6bit_6.c<3> ;
  wire \adder_6bit_6.c<4> ;
  wire \adder_6bit_6.c<5> ;
  wire \adder_6bit_6.s<0> ;
  wire \adder_6bit_6.s<1> ;
  wire \adder_6bit_6.s<2> ;
  wire \adder_6bit_6.s<3> ;
  wire \adder_6bit_6.s<4> ;
  wire \adder_6bit_6.s<5> ;
  wire \adder_6bit_6.s<6> ;
  wire \adder_6bit_6.sign ;
  wire \adder_6bit_7.a<0> ;
  wire \adder_6bit_7.a<1> ;
  wire \adder_6bit_7.a<2> ;
  wire \adder_6bit_7.a<3> ;
  wire \adder_6bit_7.a<4> ;
  wire \adder_6bit_7.a<5> ;
  wire \adder_6bit_7.b<0> ;
  wire \adder_6bit_7.b<1> ;
  wire \adder_6bit_7.b<2> ;
  wire \adder_6bit_7.b<3> ;
  wire \adder_6bit_7.b<4> ;
  wire \adder_6bit_7.b<5> ;
  wire \adder_6bit_7.c<0> ;
  wire \adder_6bit_7.c<1> ;
  wire \adder_6bit_7.c<2> ;
  wire \adder_6bit_7.c<3> ;
  wire \adder_6bit_7.c<4> ;
  wire \adder_6bit_7.c<5> ;
  wire \adder_6bit_7.s<0> ;
  wire \adder_6bit_7.s<1> ;
  wire \adder_6bit_7.s<2> ;
  wire \adder_6bit_7.s<3> ;
  wire \adder_6bit_7.s<4> ;
  wire \adder_6bit_7.s<5> ;
  wire \adder_6bit_7.s<6> ;
  wire \adder_6bit_7.sign ;
  wire \adder_7bit_0.a<0> ;
  wire \adder_7bit_0.a<1> ;
  wire \adder_7bit_0.a<2> ;
  wire \adder_7bit_0.a<3> ;
  wire \adder_7bit_0.a<4> ;
  wire \adder_7bit_0.a<5> ;
  wire \adder_7bit_0.a<6> ;
  wire \adder_7bit_0.b<0> ;
  wire \adder_7bit_0.b<1> ;
  wire \adder_7bit_0.b<2> ;
  wire \adder_7bit_0.b<3> ;
  wire \adder_7bit_0.b<4> ;
  wire \adder_7bit_0.b<5> ;
  wire \adder_7bit_0.b<6> ;
  wire \adder_7bit_0.c<0> ;
  wire \adder_7bit_0.c<1> ;
  wire \adder_7bit_0.c<2> ;
  wire \adder_7bit_0.c<3> ;
  wire \adder_7bit_0.c<4> ;
  wire \adder_7bit_0.c<5> ;
  wire \adder_7bit_0.c<6> ;
  wire \adder_7bit_0.s<0> ;
  wire \adder_7bit_0.s<1> ;
  wire \adder_7bit_0.s<2> ;
  wire \adder_7bit_0.s<3> ;
  wire \adder_7bit_0.s<4> ;
  wire \adder_7bit_0.s<5> ;
  wire \adder_7bit_0.s<6> ;
  wire \adder_7bit_0.s<7> ;
  wire \adder_7bit_0.sign ;
  wire \adder_7bit_1.a<0> ;
  wire \adder_7bit_1.a<1> ;
  wire \adder_7bit_1.a<2> ;
  wire \adder_7bit_1.a<3> ;
  wire \adder_7bit_1.a<4> ;
  wire \adder_7bit_1.a<5> ;
  wire \adder_7bit_1.a<6> ;
  wire \adder_7bit_1.b<0> ;
  wire \adder_7bit_1.b<1> ;
  wire \adder_7bit_1.b<2> ;
  wire \adder_7bit_1.b<3> ;
  wire \adder_7bit_1.b<4> ;
  wire \adder_7bit_1.b<5> ;
  wire \adder_7bit_1.b<6> ;
  wire \adder_7bit_1.c<0> ;
  wire \adder_7bit_1.c<1> ;
  wire \adder_7bit_1.c<2> ;
  wire \adder_7bit_1.c<3> ;
  wire \adder_7bit_1.c<4> ;
  wire \adder_7bit_1.c<5> ;
  wire \adder_7bit_1.c<6> ;
  wire \adder_7bit_1.s<0> ;
  wire \adder_7bit_1.s<1> ;
  wire \adder_7bit_1.s<2> ;
  wire \adder_7bit_1.s<3> ;
  wire \adder_7bit_1.s<4> ;
  wire \adder_7bit_1.s<5> ;
  wire \adder_7bit_1.s<6> ;
  wire \adder_7bit_1.s<7> ;
  wire \adder_7bit_1.sign ;
  wire \adder_7bit_2.a<0> ;
  wire \adder_7bit_2.a<1> ;
  wire \adder_7bit_2.a<2> ;
  wire \adder_7bit_2.a<3> ;
  wire \adder_7bit_2.a<4> ;
  wire \adder_7bit_2.a<5> ;
  wire \adder_7bit_2.a<6> ;
  wire \adder_7bit_2.b<0> ;
  wire \adder_7bit_2.b<1> ;
  wire \adder_7bit_2.b<2> ;
  wire \adder_7bit_2.b<3> ;
  wire \adder_7bit_2.b<4> ;
  wire \adder_7bit_2.b<5> ;
  wire \adder_7bit_2.b<6> ;
  wire \adder_7bit_2.c<0> ;
  wire \adder_7bit_2.c<1> ;
  wire \adder_7bit_2.c<2> ;
  wire \adder_7bit_2.c<3> ;
  wire \adder_7bit_2.c<4> ;
  wire \adder_7bit_2.c<5> ;
  wire \adder_7bit_2.c<6> ;
  wire \adder_7bit_2.s<0> ;
  wire \adder_7bit_2.s<1> ;
  wire \adder_7bit_2.s<2> ;
  wire \adder_7bit_2.s<3> ;
  wire \adder_7bit_2.s<4> ;
  wire \adder_7bit_2.s<5> ;
  wire \adder_7bit_2.s<6> ;
  wire \adder_7bit_2.s<7> ;
  wire \adder_7bit_2.sign ;
  wire \adder_7bit_3.a<0> ;
  wire \adder_7bit_3.a<1> ;
  wire \adder_7bit_3.a<2> ;
  wire \adder_7bit_3.a<3> ;
  wire \adder_7bit_3.a<4> ;
  wire \adder_7bit_3.a<5> ;
  wire \adder_7bit_3.a<6> ;
  wire \adder_7bit_3.b<0> ;
  wire \adder_7bit_3.b<1> ;
  wire \adder_7bit_3.b<2> ;
  wire \adder_7bit_3.b<3> ;
  wire \adder_7bit_3.b<4> ;
  wire \adder_7bit_3.b<5> ;
  wire \adder_7bit_3.b<6> ;
  wire \adder_7bit_3.c<0> ;
  wire \adder_7bit_3.c<1> ;
  wire \adder_7bit_3.c<2> ;
  wire \adder_7bit_3.c<3> ;
  wire \adder_7bit_3.c<4> ;
  wire \adder_7bit_3.c<5> ;
  wire \adder_7bit_3.c<6> ;
  wire \adder_7bit_3.s<0> ;
  wire \adder_7bit_3.s<1> ;
  wire \adder_7bit_3.s<2> ;
  wire \adder_7bit_3.s<3> ;
  wire \adder_7bit_3.s<4> ;
  wire \adder_7bit_3.s<5> ;
  wire \adder_7bit_3.s<6> ;
  wire \adder_7bit_3.s<7> ;
  wire \adder_7bit_3.sign ;
  wire \adder_8bit_0.a<0> ;
  wire \adder_8bit_0.a<1> ;
  wire \adder_8bit_0.a<2> ;
  wire \adder_8bit_0.a<3> ;
  wire \adder_8bit_0.a<4> ;
  wire \adder_8bit_0.a<5> ;
  wire \adder_8bit_0.a<6> ;
  wire \adder_8bit_0.a<7> ;
  wire \adder_8bit_0.b<0> ;
  wire \adder_8bit_0.b<1> ;
  wire \adder_8bit_0.b<2> ;
  wire \adder_8bit_0.b<3> ;
  wire \adder_8bit_0.b<4> ;
  wire \adder_8bit_0.b<5> ;
  wire \adder_8bit_0.b<6> ;
  wire \adder_8bit_0.b<7> ;
  wire \adder_8bit_0.c<0> ;
  wire \adder_8bit_0.c<1> ;
  wire \adder_8bit_0.c<2> ;
  wire \adder_8bit_0.c<3> ;
  wire \adder_8bit_0.c<4> ;
  wire \adder_8bit_0.c<5> ;
  wire \adder_8bit_0.c<6> ;
  wire \adder_8bit_0.c<7> ;
  wire \adder_8bit_0.s<0> ;
  wire \adder_8bit_0.s<1> ;
  wire \adder_8bit_0.s<2> ;
  wire \adder_8bit_0.s<3> ;
  wire \adder_8bit_0.s<4> ;
  wire \adder_8bit_0.s<5> ;
  wire \adder_8bit_0.s<6> ;
  wire \adder_8bit_0.s<7> ;
  wire \adder_8bit_0.s<8> ;
  wire \adder_8bit_0.sign ;
  wire \adder_8bit_1.a<0> ;
  wire \adder_8bit_1.a<1> ;
  wire \adder_8bit_1.a<2> ;
  wire \adder_8bit_1.a<3> ;
  wire \adder_8bit_1.a<4> ;
  wire \adder_8bit_1.a<5> ;
  wire \adder_8bit_1.a<6> ;
  wire \adder_8bit_1.a<7> ;
  wire \adder_8bit_1.b<0> ;
  wire \adder_8bit_1.b<1> ;
  wire \adder_8bit_1.b<2> ;
  wire \adder_8bit_1.b<3> ;
  wire \adder_8bit_1.b<4> ;
  wire \adder_8bit_1.b<5> ;
  wire \adder_8bit_1.b<6> ;
  wire \adder_8bit_1.b<7> ;
  wire \adder_8bit_1.c<0> ;
  wire \adder_8bit_1.c<1> ;
  wire \adder_8bit_1.c<2> ;
  wire \adder_8bit_1.c<3> ;
  wire \adder_8bit_1.c<4> ;
  wire \adder_8bit_1.c<5> ;
  wire \adder_8bit_1.c<6> ;
  wire \adder_8bit_1.c<7> ;
  wire \adder_8bit_1.s<0> ;
  wire \adder_8bit_1.s<1> ;
  wire \adder_8bit_1.s<2> ;
  wire \adder_8bit_1.s<3> ;
  wire \adder_8bit_1.s<4> ;
  wire \adder_8bit_1.s<5> ;
  wire \adder_8bit_1.s<6> ;
  wire \adder_8bit_1.s<7> ;
  wire \adder_8bit_1.s<8> ;
  wire \adder_8bit_1.sign ;
  wire \adder_9bit.a<0> ;
  wire \adder_9bit.a<1> ;
  wire \adder_9bit.a<2> ;
  wire \adder_9bit.a<3> ;
  wire \adder_9bit.a<4> ;
  wire \adder_9bit.a<5> ;
  wire \adder_9bit.a<6> ;
  wire \adder_9bit.a<7> ;
  wire \adder_9bit.a<8> ;
  wire \adder_9bit.b<0> ;
  wire \adder_9bit.b<1> ;
  wire \adder_9bit.b<2> ;
  wire \adder_9bit.b<3> ;
  wire \adder_9bit.b<4> ;
  wire \adder_9bit.b<5> ;
  wire \adder_9bit.b<6> ;
  wire \adder_9bit.b<7> ;
  wire \adder_9bit.b<8> ;
  wire \adder_9bit.c<0> ;
  wire \adder_9bit.c<1> ;
  wire \adder_9bit.c<2> ;
  wire \adder_9bit.c<3> ;
  wire \adder_9bit.c<4> ;
  wire \adder_9bit.c<5> ;
  wire \adder_9bit.c<6> ;
  wire \adder_9bit.c<7> ;
  wire \adder_9bit.c<8> ;
  wire \adder_9bit.s<0> ;
  wire \adder_9bit.s<1> ;
  wire \adder_9bit.s<2> ;
  wire \adder_9bit.s<3> ;
  wire \adder_9bit.s<4> ;
  wire \adder_9bit.s<5> ;
  wire \adder_9bit.s<6> ;
  wire \adder_9bit.s<7> ;
  wire \adder_9bit.s<8> ;
  wire \adder_9bit.s<9> ;
  wire \adder_9bit.sign ;
  input \in_0<0> ;
  input \in_0<1> ;
  input \in_0<2> ;
  input \in_0<3> ;
  input \in_10<0> ;
  input \in_10<1> ;
  input \in_10<2> ;
  input \in_10<3> ;
  input \in_11<0> ;
  input \in_11<1> ;
  input \in_11<2> ;
  input \in_11<3> ;
  input \in_12<0> ;
  input \in_12<1> ;
  input \in_12<2> ;
  input \in_12<3> ;
  input \in_13<0> ;
  input \in_13<1> ;
  input \in_13<2> ;
  input \in_13<3> ;
  input \in_14<0> ;
  input \in_14<1> ;
  input \in_14<2> ;
  input \in_14<3> ;
  input \in_15<0> ;
  input \in_15<1> ;
  input \in_15<2> ;
  input \in_15<3> ;
  input \in_16<0> ;
  input \in_16<1> ;
  input \in_16<2> ;
  input \in_16<3> ;
  input \in_17<0> ;
  input \in_17<1> ;
  input \in_17<2> ;
  input \in_17<3> ;
  input \in_18<0> ;
  input \in_18<1> ;
  input \in_18<2> ;
  input \in_18<3> ;
  input \in_19<0> ;
  input \in_19<1> ;
  input \in_19<2> ;
  input \in_19<3> ;
  input \in_1<0> ;
  input \in_1<1> ;
  input \in_1<2> ;
  input \in_1<3> ;
  input \in_20<0> ;
  input \in_20<1> ;
  input \in_20<2> ;
  input \in_20<3> ;
  input \in_21<0> ;
  input \in_21<1> ;
  input \in_21<2> ;
  input \in_21<3> ;
  input \in_22<0> ;
  input \in_22<1> ;
  input \in_22<2> ;
  input \in_22<3> ;
  input \in_23<0> ;
  input \in_23<1> ;
  input \in_23<2> ;
  input \in_23<3> ;
  input \in_24<0> ;
  input \in_24<1> ;
  input \in_24<2> ;
  input \in_24<3> ;
  input \in_25<0> ;
  input \in_25<1> ;
  input \in_25<2> ;
  input \in_25<3> ;
  input \in_26<0> ;
  input \in_26<1> ;
  input \in_26<2> ;
  input \in_26<3> ;
  input \in_27<0> ;
  input \in_27<1> ;
  input \in_27<2> ;
  input \in_27<3> ;
  input \in_28<0> ;
  input \in_28<1> ;
  input \in_28<2> ;
  input \in_28<3> ;
  input \in_29<0> ;
  input \in_29<1> ;
  input \in_29<2> ;
  input \in_29<3> ;
  input \in_2<0> ;
  input \in_2<1> ;
  input \in_2<2> ;
  input \in_2<3> ;
  input \in_30<0> ;
  input \in_30<1> ;
  input \in_30<2> ;
  input \in_30<3> ;
  input \in_31<0> ;
  input \in_31<1> ;
  input \in_31<2> ;
  input \in_31<3> ;
  input \in_32<0> ;
  input \in_32<1> ;
  input \in_32<2> ;
  input \in_32<3> ;
  input \in_33<0> ;
  input \in_33<1> ;
  input \in_33<2> ;
  input \in_33<3> ;
  input \in_34<0> ;
  input \in_34<1> ;
  input \in_34<2> ;
  input \in_34<3> ;
  input \in_35<0> ;
  input \in_35<1> ;
  input \in_35<2> ;
  input \in_35<3> ;
  input \in_36<0> ;
  input \in_36<1> ;
  input \in_36<2> ;
  input \in_36<3> ;
  input \in_37<0> ;
  input \in_37<1> ;
  input \in_37<2> ;
  input \in_37<3> ;
  input \in_38<0> ;
  input \in_38<1> ;
  input \in_38<2> ;
  input \in_38<3> ;
  input \in_39<0> ;
  input \in_39<1> ;
  input \in_39<2> ;
  input \in_39<3> ;
  input \in_3<0> ;
  input \in_3<1> ;
  input \in_3<2> ;
  input \in_3<3> ;
  input \in_40<0> ;
  input \in_40<1> ;
  input \in_40<2> ;
  input \in_40<3> ;
  input \in_41<0> ;
  input \in_41<1> ;
  input \in_41<2> ;
  input \in_41<3> ;
  input \in_42<0> ;
  input \in_42<1> ;
  input \in_42<2> ;
  input \in_42<3> ;
  input \in_43<0> ;
  input \in_43<1> ;
  input \in_43<2> ;
  input \in_43<3> ;
  input \in_44<0> ;
  input \in_44<1> ;
  input \in_44<2> ;
  input \in_44<3> ;
  input \in_45<0> ;
  input \in_45<1> ;
  input \in_45<2> ;
  input \in_45<3> ;
  input \in_46<0> ;
  input \in_46<1> ;
  input \in_46<2> ;
  input \in_46<3> ;
  input \in_47<0> ;
  input \in_47<1> ;
  input \in_47<2> ;
  input \in_47<3> ;
  input \in_48<0> ;
  input \in_48<1> ;
  input \in_48<2> ;
  input \in_48<3> ;
  input \in_49<0> ;
  input \in_49<1> ;
  input \in_49<2> ;
  input \in_49<3> ;
  input \in_4<0> ;
  input \in_4<1> ;
  input \in_4<2> ;
  input \in_4<3> ;
  input \in_50<0> ;
  input \in_50<1> ;
  input \in_50<2> ;
  input \in_50<3> ;
  input \in_51<0> ;
  input \in_51<1> ;
  input \in_51<2> ;
  input \in_51<3> ;
  input \in_52<0> ;
  input \in_52<1> ;
  input \in_52<2> ;
  input \in_52<3> ;
  input \in_53<0> ;
  input \in_53<1> ;
  input \in_53<2> ;
  input \in_53<3> ;
  input \in_54<0> ;
  input \in_54<1> ;
  input \in_54<2> ;
  input \in_54<3> ;
  input \in_55<0> ;
  input \in_55<1> ;
  input \in_55<2> ;
  input \in_55<3> ;
  input \in_56<0> ;
  input \in_56<1> ;
  input \in_56<2> ;
  input \in_56<3> ;
  input \in_57<0> ;
  input \in_57<1> ;
  input \in_57<2> ;
  input \in_57<3> ;
  input \in_58<0> ;
  input \in_58<1> ;
  input \in_58<2> ;
  input \in_58<3> ;
  input \in_59<0> ;
  input \in_59<1> ;
  input \in_59<2> ;
  input \in_59<3> ;
  input \in_5<0> ;
  input \in_5<1> ;
  input \in_5<2> ;
  input \in_5<3> ;
  input \in_60<0> ;
  input \in_60<1> ;
  input \in_60<2> ;
  input \in_60<3> ;
  input \in_61<0> ;
  input \in_61<1> ;
  input \in_61<2> ;
  input \in_61<3> ;
  input \in_62<0> ;
  input \in_62<1> ;
  input \in_62<2> ;
  input \in_62<3> ;
  input \in_63<0> ;
  input \in_63<1> ;
  input \in_63<2> ;
  input \in_63<3> ;
  input \in_6<0> ;
  input \in_6<1> ;
  input \in_6<2> ;
  input \in_6<3> ;
  input \in_7<0> ;
  input \in_7<1> ;
  input \in_7<2> ;
  input \in_7<3> ;
  input \in_8<0> ;
  input \in_8<1> ;
  input \in_8<2> ;
  input \in_8<3> ;
  input \in_9<0> ;
  input \in_9<1> ;
  input \in_9<2> ;
  input \in_9<3> ;
  output \out<0> ;
  output \out<1> ;
  output \out<2> ;
  output \out<3> ;
  output \out<4> ;
  output \out<5> ;
  output \out<6> ;
  output \out<7> ;
  output \out<8> ;
  output \out<9> ;
  input sign_weight;
  wire \sum_4bit_0<0> ;
  wire \sum_4bit_0<1> ;
  wire \sum_4bit_0<2> ;
  wire \sum_4bit_0<3> ;
  wire \sum_4bit_0<4> ;
  wire \sum_4bit_10<0> ;
  wire \sum_4bit_10<1> ;
  wire \sum_4bit_10<2> ;
  wire \sum_4bit_10<3> ;
  wire \sum_4bit_10<4> ;
  wire \sum_4bit_11<0> ;
  wire \sum_4bit_11<1> ;
  wire \sum_4bit_11<2> ;
  wire \sum_4bit_11<3> ;
  wire \sum_4bit_11<4> ;
  wire \sum_4bit_12<0> ;
  wire \sum_4bit_12<1> ;
  wire \sum_4bit_12<2> ;
  wire \sum_4bit_12<3> ;
  wire \sum_4bit_12<4> ;
  wire \sum_4bit_13<0> ;
  wire \sum_4bit_13<1> ;
  wire \sum_4bit_13<2> ;
  wire \sum_4bit_13<3> ;
  wire \sum_4bit_13<4> ;
  wire \sum_4bit_14<0> ;
  wire \sum_4bit_14<1> ;
  wire \sum_4bit_14<2> ;
  wire \sum_4bit_14<3> ;
  wire \sum_4bit_14<4> ;
  wire \sum_4bit_15<0> ;
  wire \sum_4bit_15<1> ;
  wire \sum_4bit_15<2> ;
  wire \sum_4bit_15<3> ;
  wire \sum_4bit_15<4> ;
  wire \sum_4bit_16<0> ;
  wire \sum_4bit_16<1> ;
  wire \sum_4bit_16<2> ;
  wire \sum_4bit_16<3> ;
  wire \sum_4bit_16<4> ;
  wire \sum_4bit_17<0> ;
  wire \sum_4bit_17<1> ;
  wire \sum_4bit_17<2> ;
  wire \sum_4bit_17<3> ;
  wire \sum_4bit_17<4> ;
  wire \sum_4bit_18<0> ;
  wire \sum_4bit_18<1> ;
  wire \sum_4bit_18<2> ;
  wire \sum_4bit_18<3> ;
  wire \sum_4bit_18<4> ;
  wire \sum_4bit_19<0> ;
  wire \sum_4bit_19<1> ;
  wire \sum_4bit_19<2> ;
  wire \sum_4bit_19<3> ;
  wire \sum_4bit_19<4> ;
  wire \sum_4bit_1<0> ;
  wire \sum_4bit_1<1> ;
  wire \sum_4bit_1<2> ;
  wire \sum_4bit_1<3> ;
  wire \sum_4bit_1<4> ;
  wire \sum_4bit_20<0> ;
  wire \sum_4bit_20<1> ;
  wire \sum_4bit_20<2> ;
  wire \sum_4bit_20<3> ;
  wire \sum_4bit_20<4> ;
  wire \sum_4bit_21<0> ;
  wire \sum_4bit_21<1> ;
  wire \sum_4bit_21<2> ;
  wire \sum_4bit_21<3> ;
  wire \sum_4bit_21<4> ;
  wire \sum_4bit_22<0> ;
  wire \sum_4bit_22<1> ;
  wire \sum_4bit_22<2> ;
  wire \sum_4bit_22<3> ;
  wire \sum_4bit_22<4> ;
  wire \sum_4bit_23<0> ;
  wire \sum_4bit_23<1> ;
  wire \sum_4bit_23<2> ;
  wire \sum_4bit_23<3> ;
  wire \sum_4bit_23<4> ;
  wire \sum_4bit_24<0> ;
  wire \sum_4bit_24<1> ;
  wire \sum_4bit_24<2> ;
  wire \sum_4bit_24<3> ;
  wire \sum_4bit_24<4> ;
  wire \sum_4bit_25<0> ;
  wire \sum_4bit_25<1> ;
  wire \sum_4bit_25<2> ;
  wire \sum_4bit_25<3> ;
  wire \sum_4bit_25<4> ;
  wire \sum_4bit_26<0> ;
  wire \sum_4bit_26<1> ;
  wire \sum_4bit_26<2> ;
  wire \sum_4bit_26<3> ;
  wire \sum_4bit_26<4> ;
  wire \sum_4bit_27<0> ;
  wire \sum_4bit_27<1> ;
  wire \sum_4bit_27<2> ;
  wire \sum_4bit_27<3> ;
  wire \sum_4bit_27<4> ;
  wire \sum_4bit_28<0> ;
  wire \sum_4bit_28<1> ;
  wire \sum_4bit_28<2> ;
  wire \sum_4bit_28<3> ;
  wire \sum_4bit_28<4> ;
  wire \sum_4bit_29<0> ;
  wire \sum_4bit_29<1> ;
  wire \sum_4bit_29<2> ;
  wire \sum_4bit_29<3> ;
  wire \sum_4bit_29<4> ;
  wire \sum_4bit_2<0> ;
  wire \sum_4bit_2<1> ;
  wire \sum_4bit_2<2> ;
  wire \sum_4bit_2<3> ;
  wire \sum_4bit_2<4> ;
  wire \sum_4bit_30<0> ;
  wire \sum_4bit_30<1> ;
  wire \sum_4bit_30<2> ;
  wire \sum_4bit_30<3> ;
  wire \sum_4bit_30<4> ;
  wire \sum_4bit_31<0> ;
  wire \sum_4bit_31<1> ;
  wire \sum_4bit_31<2> ;
  wire \sum_4bit_31<3> ;
  wire \sum_4bit_31<4> ;
  wire \sum_4bit_3<0> ;
  wire \sum_4bit_3<1> ;
  wire \sum_4bit_3<2> ;
  wire \sum_4bit_3<3> ;
  wire \sum_4bit_3<4> ;
  wire \sum_4bit_4<0> ;
  wire \sum_4bit_4<1> ;
  wire \sum_4bit_4<2> ;
  wire \sum_4bit_4<3> ;
  wire \sum_4bit_4<4> ;
  wire \sum_4bit_5<0> ;
  wire \sum_4bit_5<1> ;
  wire \sum_4bit_5<2> ;
  wire \sum_4bit_5<3> ;
  wire \sum_4bit_5<4> ;
  wire \sum_4bit_6<0> ;
  wire \sum_4bit_6<1> ;
  wire \sum_4bit_6<2> ;
  wire \sum_4bit_6<3> ;
  wire \sum_4bit_6<4> ;
  wire \sum_4bit_7<0> ;
  wire \sum_4bit_7<1> ;
  wire \sum_4bit_7<2> ;
  wire \sum_4bit_7<3> ;
  wire \sum_4bit_7<4> ;
  wire \sum_4bit_8<0> ;
  wire \sum_4bit_8<1> ;
  wire \sum_4bit_8<2> ;
  wire \sum_4bit_8<3> ;
  wire \sum_4bit_8<4> ;
  wire \sum_4bit_9<0> ;
  wire \sum_4bit_9<1> ;
  wire \sum_4bit_9<2> ;
  wire \sum_4bit_9<3> ;
  wire \sum_4bit_9<4> ;
  wire \sum_5bit_0<0> ;
  wire \sum_5bit_0<1> ;
  wire \sum_5bit_0<2> ;
  wire \sum_5bit_0<3> ;
  wire \sum_5bit_0<4> ;
  wire \sum_5bit_0<5> ;
  wire \sum_5bit_10<0> ;
  wire \sum_5bit_10<1> ;
  wire \sum_5bit_10<2> ;
  wire \sum_5bit_10<3> ;
  wire \sum_5bit_10<4> ;
  wire \sum_5bit_10<5> ;
  wire \sum_5bit_11<0> ;
  wire \sum_5bit_11<1> ;
  wire \sum_5bit_11<2> ;
  wire \sum_5bit_11<3> ;
  wire \sum_5bit_11<4> ;
  wire \sum_5bit_11<5> ;
  wire \sum_5bit_12<0> ;
  wire \sum_5bit_12<1> ;
  wire \sum_5bit_12<2> ;
  wire \sum_5bit_12<3> ;
  wire \sum_5bit_12<4> ;
  wire \sum_5bit_12<5> ;
  wire \sum_5bit_13<0> ;
  wire \sum_5bit_13<1> ;
  wire \sum_5bit_13<2> ;
  wire \sum_5bit_13<3> ;
  wire \sum_5bit_13<4> ;
  wire \sum_5bit_13<5> ;
  wire \sum_5bit_14<0> ;
  wire \sum_5bit_14<1> ;
  wire \sum_5bit_14<2> ;
  wire \sum_5bit_14<3> ;
  wire \sum_5bit_14<4> ;
  wire \sum_5bit_14<5> ;
  wire \sum_5bit_15<0> ;
  wire \sum_5bit_15<1> ;
  wire \sum_5bit_15<2> ;
  wire \sum_5bit_15<3> ;
  wire \sum_5bit_15<4> ;
  wire \sum_5bit_15<5> ;
  wire \sum_5bit_1<0> ;
  wire \sum_5bit_1<1> ;
  wire \sum_5bit_1<2> ;
  wire \sum_5bit_1<3> ;
  wire \sum_5bit_1<4> ;
  wire \sum_5bit_1<5> ;
  wire \sum_5bit_2<0> ;
  wire \sum_5bit_2<1> ;
  wire \sum_5bit_2<2> ;
  wire \sum_5bit_2<3> ;
  wire \sum_5bit_2<4> ;
  wire \sum_5bit_2<5> ;
  wire \sum_5bit_3<0> ;
  wire \sum_5bit_3<1> ;
  wire \sum_5bit_3<2> ;
  wire \sum_5bit_3<3> ;
  wire \sum_5bit_3<4> ;
  wire \sum_5bit_3<5> ;
  wire \sum_5bit_4<0> ;
  wire \sum_5bit_4<1> ;
  wire \sum_5bit_4<2> ;
  wire \sum_5bit_4<3> ;
  wire \sum_5bit_4<4> ;
  wire \sum_5bit_4<5> ;
  wire \sum_5bit_5<0> ;
  wire \sum_5bit_5<1> ;
  wire \sum_5bit_5<2> ;
  wire \sum_5bit_5<3> ;
  wire \sum_5bit_5<4> ;
  wire \sum_5bit_5<5> ;
  wire \sum_5bit_6<0> ;
  wire \sum_5bit_6<1> ;
  wire \sum_5bit_6<2> ;
  wire \sum_5bit_6<3> ;
  wire \sum_5bit_6<4> ;
  wire \sum_5bit_6<5> ;
  wire \sum_5bit_7<0> ;
  wire \sum_5bit_7<1> ;
  wire \sum_5bit_7<2> ;
  wire \sum_5bit_7<3> ;
  wire \sum_5bit_7<4> ;
  wire \sum_5bit_7<5> ;
  wire \sum_5bit_8<0> ;
  wire \sum_5bit_8<1> ;
  wire \sum_5bit_8<2> ;
  wire \sum_5bit_8<3> ;
  wire \sum_5bit_8<4> ;
  wire \sum_5bit_8<5> ;
  wire \sum_5bit_9<0> ;
  wire \sum_5bit_9<1> ;
  wire \sum_5bit_9<2> ;
  wire \sum_5bit_9<3> ;
  wire \sum_5bit_9<4> ;
  wire \sum_5bit_9<5> ;
  wire \sum_6bit_0<0> ;
  wire \sum_6bit_0<1> ;
  wire \sum_6bit_0<2> ;
  wire \sum_6bit_0<3> ;
  wire \sum_6bit_0<4> ;
  wire \sum_6bit_0<5> ;
  wire \sum_6bit_0<6> ;
  wire \sum_6bit_1<0> ;
  wire \sum_6bit_1<1> ;
  wire \sum_6bit_1<2> ;
  wire \sum_6bit_1<3> ;
  wire \sum_6bit_1<4> ;
  wire \sum_6bit_1<5> ;
  wire \sum_6bit_1<6> ;
  wire \sum_6bit_2<0> ;
  wire \sum_6bit_2<1> ;
  wire \sum_6bit_2<2> ;
  wire \sum_6bit_2<3> ;
  wire \sum_6bit_2<4> ;
  wire \sum_6bit_2<5> ;
  wire \sum_6bit_2<6> ;
  wire \sum_6bit_3<0> ;
  wire \sum_6bit_3<1> ;
  wire \sum_6bit_3<2> ;
  wire \sum_6bit_3<3> ;
  wire \sum_6bit_3<4> ;
  wire \sum_6bit_3<5> ;
  wire \sum_6bit_3<6> ;
  wire \sum_6bit_4<0> ;
  wire \sum_6bit_4<1> ;
  wire \sum_6bit_4<2> ;
  wire \sum_6bit_4<3> ;
  wire \sum_6bit_4<4> ;
  wire \sum_6bit_4<5> ;
  wire \sum_6bit_4<6> ;
  wire \sum_6bit_5<0> ;
  wire \sum_6bit_5<1> ;
  wire \sum_6bit_5<2> ;
  wire \sum_6bit_5<3> ;
  wire \sum_6bit_5<4> ;
  wire \sum_6bit_5<5> ;
  wire \sum_6bit_5<6> ;
  wire \sum_6bit_6<0> ;
  wire \sum_6bit_6<1> ;
  wire \sum_6bit_6<2> ;
  wire \sum_6bit_6<3> ;
  wire \sum_6bit_6<4> ;
  wire \sum_6bit_6<5> ;
  wire \sum_6bit_6<6> ;
  wire \sum_6bit_7<0> ;
  wire \sum_6bit_7<1> ;
  wire \sum_6bit_7<2> ;
  wire \sum_6bit_7<3> ;
  wire \sum_6bit_7<4> ;
  wire \sum_6bit_7<5> ;
  wire \sum_6bit_7<6> ;
  wire \sum_7bit_0<0> ;
  wire \sum_7bit_0<1> ;
  wire \sum_7bit_0<2> ;
  wire \sum_7bit_0<3> ;
  wire \sum_7bit_0<4> ;
  wire \sum_7bit_0<5> ;
  wire \sum_7bit_0<6> ;
  wire \sum_7bit_0<7> ;
  wire \sum_7bit_1<0> ;
  wire \sum_7bit_1<1> ;
  wire \sum_7bit_1<2> ;
  wire \sum_7bit_1<3> ;
  wire \sum_7bit_1<4> ;
  wire \sum_7bit_1<5> ;
  wire \sum_7bit_1<6> ;
  wire \sum_7bit_1<7> ;
  wire \sum_7bit_2<0> ;
  wire \sum_7bit_2<1> ;
  wire \sum_7bit_2<2> ;
  wire \sum_7bit_2<3> ;
  wire \sum_7bit_2<4> ;
  wire \sum_7bit_2<5> ;
  wire \sum_7bit_2<6> ;
  wire \sum_7bit_2<7> ;
  wire \sum_7bit_3<0> ;
  wire \sum_7bit_3<1> ;
  wire \sum_7bit_3<2> ;
  wire \sum_7bit_3<3> ;
  wire \sum_7bit_3<4> ;
  wire \sum_7bit_3<5> ;
  wire \sum_7bit_3<6> ;
  wire \sum_7bit_3<7> ;
  wire \sum_8bit_0<0> ;
  wire \sum_8bit_0<1> ;
  wire \sum_8bit_0<2> ;
  wire \sum_8bit_0<3> ;
  wire \sum_8bit_0<4> ;
  wire \sum_8bit_0<5> ;
  wire \sum_8bit_0<6> ;
  wire \sum_8bit_0<7> ;
  wire \sum_8bit_0<8> ;
  wire \sum_8bit_1<0> ;
  wire \sum_8bit_1<1> ;
  wire \sum_8bit_1<2> ;
  wire \sum_8bit_1<3> ;
  wire \sum_8bit_1<4> ;
  wire \sum_8bit_1<5> ;
  wire \sum_8bit_1<6> ;
  wire \sum_8bit_1<7> ;
  wire \sum_8bit_1<8> ;
  full_adder \adder_4bit_0.fa_1  (    .a(\in_0<1> ),    .b(\in_1<1> ),    .cin(\adder_4bit_0.c<0> ),    .cout(\adder_4bit_0.c<1> ),    .s(\adder_4bit_0.s<1> )
  );
  full_adder \adder_4bit_0.fa_2  (    .a(\in_0<2> ),    .b(\in_1<2> ),    .cin(\adder_4bit_0.c<1> ),    .cout(\adder_4bit_0.c<2> ),    .s(\adder_4bit_0.s<2> )
  );
  full_adder \adder_4bit_0.fa_3  (    .a(\in_0<3> ),    .b(\in_1<3> ),    .cin(\adder_4bit_0.c<2> ),    .cout(\adder_4bit_0.c<3> ),    .s(\adder_4bit_0.s<3> )
  );
  adder_sign_extension \adder_4bit_0.fa_4  (    .a(\in_0<3> ),    .b(\in_1<3> ),    .cin(\adder_4bit_0.c<3> ),    .s(\adder_4bit_0.s<4> ),    .sign(sign_weight)
  );
  half_adder \adder_4bit_0.ha_0  (    .a(\in_0<0> ),    .b(\in_1<0> ),    .cout(\adder_4bit_0.c<0> ),    .s(\adder_4bit_0.s<0> )
  );
  full_adder \adder_4bit_1.fa_1  (    .a(\in_2<1> ),    .b(\in_3<1> ),    .cin(\adder_4bit_1.c<0> ),    .cout(\adder_4bit_1.c<1> ),    .s(\adder_4bit_1.s<1> )
  );
  full_adder \adder_4bit_1.fa_2  (    .a(\in_2<2> ),    .b(\in_3<2> ),    .cin(\adder_4bit_1.c<1> ),    .cout(\adder_4bit_1.c<2> ),    .s(\adder_4bit_1.s<2> )
  );
  full_adder \adder_4bit_1.fa_3  (    .a(\in_2<3> ),    .b(\in_3<3> ),    .cin(\adder_4bit_1.c<2> ),    .cout(\adder_4bit_1.c<3> ),    .s(\adder_4bit_1.s<3> )
  );
  adder_sign_extension \adder_4bit_1.fa_4  (    .a(\in_2<3> ),    .b(\in_3<3> ),    .cin(\adder_4bit_1.c<3> ),    .s(\adder_4bit_1.s<4> ),    .sign(sign_weight)
  );
  half_adder \adder_4bit_1.ha_0  (    .a(\in_2<0> ),    .b(\in_3<0> ),    .cout(\adder_4bit_1.c<0> ),    .s(\adder_4bit_1.s<0> )
  );
  full_adder \adder_4bit_10.fa_1  (    .a(\in_20<1> ),    .b(\in_21<1> ),    .cin(\adder_4bit_10.c<0> ),    .cout(\adder_4bit_10.c<1> ),    .s(\adder_4bit_10.s<1> )
  );
  full_adder \adder_4bit_10.fa_2  (    .a(\in_20<2> ),    .b(\in_21<2> ),    .cin(\adder_4bit_10.c<1> ),    .cout(\adder_4bit_10.c<2> ),    .s(\adder_4bit_10.s<2> )
  );
  full_adder \adder_4bit_10.fa_3  (    .a(\in_20<3> ),    .b(\in_21<3> ),    .cin(\adder_4bit_10.c<2> ),    .cout(\adder_4bit_10.c<3> ),    .s(\adder_4bit_10.s<3> )
  );
  adder_sign_extension \adder_4bit_10.fa_4  (    .a(\in_20<3> ),    .b(\in_21<3> ),    .cin(\adder_4bit_10.c<3> ),    .s(\adder_4bit_10.s<4> ),    .sign(sign_weight)
  );
  half_adder \adder_4bit_10.ha_0  (    .a(\in_20<0> ),    .b(\in_21<0> ),    .cout(\adder_4bit_10.c<0> ),    .s(\adder_4bit_10.s<0> )
  );
  full_adder \adder_4bit_11.fa_1  (    .a(\in_22<1> ),    .b(\in_23<1> ),    .cin(\adder_4bit_11.c<0> ),    .cout(\adder_4bit_11.c<1> ),    .s(\adder_4bit_11.s<1> )
  );
  full_adder \adder_4bit_11.fa_2  (    .a(\in_22<2> ),    .b(\in_23<2> ),    .cin(\adder_4bit_11.c<1> ),    .cout(\adder_4bit_11.c<2> ),    .s(\adder_4bit_11.s<2> )
  );
  full_adder \adder_4bit_11.fa_3  (    .a(\in_22<3> ),    .b(\in_23<3> ),    .cin(\adder_4bit_11.c<2> ),    .cout(\adder_4bit_11.c<3> ),    .s(\adder_4bit_11.s<3> )
  );
  adder_sign_extension \adder_4bit_11.fa_4  (    .a(\in_22<3> ),    .b(\in_23<3> ),    .cin(\adder_4bit_11.c<3> ),    .s(\adder_4bit_11.s<4> ),    .sign(sign_weight)
  );
  half_adder \adder_4bit_11.ha_0  (    .a(\in_22<0> ),    .b(\in_23<0> ),    .cout(\adder_4bit_11.c<0> ),    .s(\adder_4bit_11.s<0> )
  );
  full_adder \adder_4bit_12.fa_1  (    .a(\in_24<1> ),    .b(\in_25<1> ),    .cin(\adder_4bit_12.c<0> ),    .cout(\adder_4bit_12.c<1> ),    .s(\adder_4bit_12.s<1> )
  );
  full_adder \adder_4bit_12.fa_2  (    .a(\in_24<2> ),    .b(\in_25<2> ),    .cin(\adder_4bit_12.c<1> ),    .cout(\adder_4bit_12.c<2> ),    .s(\adder_4bit_12.s<2> )
  );
  full_adder \adder_4bit_12.fa_3  (    .a(\in_24<3> ),    .b(\in_25<3> ),    .cin(\adder_4bit_12.c<2> ),    .cout(\adder_4bit_12.c<3> ),    .s(\adder_4bit_12.s<3> )
  );
  adder_sign_extension \adder_4bit_12.fa_4  (    .a(\in_24<3> ),    .b(\in_25<3> ),    .cin(\adder_4bit_12.c<3> ),    .s(\adder_4bit_12.s<4> ),    .sign(sign_weight)
  );
  half_adder \adder_4bit_12.ha_0  (    .a(\in_24<0> ),    .b(\in_25<0> ),    .cout(\adder_4bit_12.c<0> ),    .s(\adder_4bit_12.s<0> )
  );
  full_adder \adder_4bit_13.fa_1  (    .a(\in_26<1> ),    .b(\in_27<1> ),    .cin(\adder_4bit_13.c<0> ),    .cout(\adder_4bit_13.c<1> ),    .s(\adder_4bit_13.s<1> )
  );
  full_adder \adder_4bit_13.fa_2  (    .a(\in_26<2> ),    .b(\in_27<2> ),    .cin(\adder_4bit_13.c<1> ),    .cout(\adder_4bit_13.c<2> ),    .s(\adder_4bit_13.s<2> )
  );
  full_adder \adder_4bit_13.fa_3  (    .a(\in_26<3> ),    .b(\in_27<3> ),    .cin(\adder_4bit_13.c<2> ),    .cout(\adder_4bit_13.c<3> ),    .s(\adder_4bit_13.s<3> )
  );
  adder_sign_extension \adder_4bit_13.fa_4  (    .a(\in_26<3> ),    .b(\in_27<3> ),    .cin(\adder_4bit_13.c<3> ),    .s(\adder_4bit_13.s<4> ),    .sign(sign_weight)
  );
  half_adder \adder_4bit_13.ha_0  (    .a(\in_26<0> ),    .b(\in_27<0> ),    .cout(\adder_4bit_13.c<0> ),    .s(\adder_4bit_13.s<0> )
  );
  full_adder \adder_4bit_14.fa_1  (    .a(\in_28<1> ),    .b(\in_29<1> ),    .cin(\adder_4bit_14.c<0> ),    .cout(\adder_4bit_14.c<1> ),    .s(\adder_4bit_14.s<1> )
  );
  full_adder \adder_4bit_14.fa_2  (    .a(\in_28<2> ),    .b(\in_29<2> ),    .cin(\adder_4bit_14.c<1> ),    .cout(\adder_4bit_14.c<2> ),    .s(\adder_4bit_14.s<2> )
  );
  full_adder \adder_4bit_14.fa_3  (    .a(\in_28<3> ),    .b(\in_29<3> ),    .cin(\adder_4bit_14.c<2> ),    .cout(\adder_4bit_14.c<3> ),    .s(\adder_4bit_14.s<3> )
  );
  adder_sign_extension \adder_4bit_14.fa_4  (    .a(\in_28<3> ),    .b(\in_29<3> ),    .cin(\adder_4bit_14.c<3> ),    .s(\adder_4bit_14.s<4> ),    .sign(sign_weight)
  );
  half_adder \adder_4bit_14.ha_0  (    .a(\in_28<0> ),    .b(\in_29<0> ),    .cout(\adder_4bit_14.c<0> ),    .s(\adder_4bit_14.s<0> )
  );
  full_adder \adder_4bit_15.fa_1  (    .a(\in_30<1> ),    .b(\in_31<1> ),    .cin(\adder_4bit_15.c<0> ),    .cout(\adder_4bit_15.c<1> ),    .s(\adder_4bit_15.s<1> )
  );
  full_adder \adder_4bit_15.fa_2  (    .a(\in_30<2> ),    .b(\in_31<2> ),    .cin(\adder_4bit_15.c<1> ),    .cout(\adder_4bit_15.c<2> ),    .s(\adder_4bit_15.s<2> )
  );
  full_adder \adder_4bit_15.fa_3  (    .a(\in_30<3> ),    .b(\in_31<3> ),    .cin(\adder_4bit_15.c<2> ),    .cout(\adder_4bit_15.c<3> ),    .s(\adder_4bit_15.s<3> )
  );
  adder_sign_extension \adder_4bit_15.fa_4  (    .a(\in_30<3> ),    .b(\in_31<3> ),    .cin(\adder_4bit_15.c<3> ),    .s(\adder_4bit_15.s<4> ),    .sign(sign_weight)
  );
  half_adder \adder_4bit_15.ha_0  (    .a(\in_30<0> ),    .b(\in_31<0> ),    .cout(\adder_4bit_15.c<0> ),    .s(\adder_4bit_15.s<0> )
  );
  full_adder \adder_4bit_16.fa_1  (    .a(\in_32<1> ),    .b(\in_33<1> ),    .cin(\adder_4bit_16.c<0> ),    .cout(\adder_4bit_16.c<1> ),    .s(\adder_4bit_16.s<1> )
  );
  full_adder \adder_4bit_16.fa_2  (    .a(\in_32<2> ),    .b(\in_33<2> ),    .cin(\adder_4bit_16.c<1> ),    .cout(\adder_4bit_16.c<2> ),    .s(\adder_4bit_16.s<2> )
  );
  full_adder \adder_4bit_16.fa_3  (    .a(\in_32<3> ),    .b(\in_33<3> ),    .cin(\adder_4bit_16.c<2> ),    .cout(\adder_4bit_16.c<3> ),    .s(\adder_4bit_16.s<3> )
  );
  adder_sign_extension \adder_4bit_16.fa_4  (    .a(\in_32<3> ),    .b(\in_33<3> ),    .cin(\adder_4bit_16.c<3> ),    .s(\adder_4bit_16.s<4> ),    .sign(sign_weight)
  );
  half_adder \adder_4bit_16.ha_0  (    .a(\in_32<0> ),    .b(\in_33<0> ),    .cout(\adder_4bit_16.c<0> ),    .s(\adder_4bit_16.s<0> )
  );
  full_adder \adder_4bit_17.fa_1  (    .a(\in_34<1> ),    .b(\in_35<1> ),    .cin(\adder_4bit_17.c<0> ),    .cout(\adder_4bit_17.c<1> ),    .s(\adder_4bit_17.s<1> )
  );
  full_adder \adder_4bit_17.fa_2  (    .a(\in_34<2> ),    .b(\in_35<2> ),    .cin(\adder_4bit_17.c<1> ),    .cout(\adder_4bit_17.c<2> ),    .s(\adder_4bit_17.s<2> )
  );
  full_adder \adder_4bit_17.fa_3  (    .a(\in_34<3> ),    .b(\in_35<3> ),    .cin(\adder_4bit_17.c<2> ),    .cout(\adder_4bit_17.c<3> ),    .s(\adder_4bit_17.s<3> )
  );
  adder_sign_extension \adder_4bit_17.fa_4  (    .a(\in_34<3> ),    .b(\in_35<3> ),    .cin(\adder_4bit_17.c<3> ),    .s(\adder_4bit_17.s<4> ),    .sign(sign_weight)
  );
  half_adder \adder_4bit_17.ha_0  (    .a(\in_34<0> ),    .b(\in_35<0> ),    .cout(\adder_4bit_17.c<0> ),    .s(\adder_4bit_17.s<0> )
  );
  full_adder \adder_4bit_18.fa_1  (    .a(\in_36<1> ),    .b(\in_37<1> ),    .cin(\adder_4bit_18.c<0> ),    .cout(\adder_4bit_18.c<1> ),    .s(\adder_4bit_18.s<1> )
  );
  full_adder \adder_4bit_18.fa_2  (    .a(\in_36<2> ),    .b(\in_37<2> ),    .cin(\adder_4bit_18.c<1> ),    .cout(\adder_4bit_18.c<2> ),    .s(\adder_4bit_18.s<2> )
  );
  full_adder \adder_4bit_18.fa_3  (    .a(\in_36<3> ),    .b(\in_37<3> ),    .cin(\adder_4bit_18.c<2> ),    .cout(\adder_4bit_18.c<3> ),    .s(\adder_4bit_18.s<3> )
  );
  adder_sign_extension \adder_4bit_18.fa_4  (    .a(\in_36<3> ),    .b(\in_37<3> ),    .cin(\adder_4bit_18.c<3> ),    .s(\adder_4bit_18.s<4> ),    .sign(sign_weight)
  );
  half_adder \adder_4bit_18.ha_0  (    .a(\in_36<0> ),    .b(\in_37<0> ),    .cout(\adder_4bit_18.c<0> ),    .s(\adder_4bit_18.s<0> )
  );
  full_adder \adder_4bit_19.fa_1  (    .a(\in_38<1> ),    .b(\in_39<1> ),    .cin(\adder_4bit_19.c<0> ),    .cout(\adder_4bit_19.c<1> ),    .s(\adder_4bit_19.s<1> )
  );
  full_adder \adder_4bit_19.fa_2  (    .a(\in_38<2> ),    .b(\in_39<2> ),    .cin(\adder_4bit_19.c<1> ),    .cout(\adder_4bit_19.c<2> ),    .s(\adder_4bit_19.s<2> )
  );
  full_adder \adder_4bit_19.fa_3  (    .a(\in_38<3> ),    .b(\in_39<3> ),    .cin(\adder_4bit_19.c<2> ),    .cout(\adder_4bit_19.c<3> ),    .s(\adder_4bit_19.s<3> )
  );
  adder_sign_extension \adder_4bit_19.fa_4  (    .a(\in_38<3> ),    .b(\in_39<3> ),    .cin(\adder_4bit_19.c<3> ),    .s(\adder_4bit_19.s<4> ),    .sign(sign_weight)
  );
  half_adder \adder_4bit_19.ha_0  (    .a(\in_38<0> ),    .b(\in_39<0> ),    .cout(\adder_4bit_19.c<0> ),    .s(\adder_4bit_19.s<0> )
  );
  full_adder \adder_4bit_2.fa_1  (    .a(\in_4<1> ),    .b(\in_5<1> ),    .cin(\adder_4bit_2.c<0> ),    .cout(\adder_4bit_2.c<1> ),    .s(\adder_4bit_2.s<1> )
  );
  full_adder \adder_4bit_2.fa_2  (    .a(\in_4<2> ),    .b(\in_5<2> ),    .cin(\adder_4bit_2.c<1> ),    .cout(\adder_4bit_2.c<2> ),    .s(\adder_4bit_2.s<2> )
  );
  full_adder \adder_4bit_2.fa_3  (    .a(\in_4<3> ),    .b(\in_5<3> ),    .cin(\adder_4bit_2.c<2> ),    .cout(\adder_4bit_2.c<3> ),    .s(\adder_4bit_2.s<3> )
  );
  adder_sign_extension \adder_4bit_2.fa_4  (    .a(\in_4<3> ),    .b(\in_5<3> ),    .cin(\adder_4bit_2.c<3> ),    .s(\adder_4bit_2.s<4> ),    .sign(sign_weight)
  );
  half_adder \adder_4bit_2.ha_0  (    .a(\in_4<0> ),    .b(\in_5<0> ),    .cout(\adder_4bit_2.c<0> ),    .s(\adder_4bit_2.s<0> )
  );
  full_adder \adder_4bit_20.fa_1  (    .a(\in_40<1> ),    .b(\in_41<1> ),    .cin(\adder_4bit_20.c<0> ),    .cout(\adder_4bit_20.c<1> ),    .s(\adder_4bit_20.s<1> )
  );
  full_adder \adder_4bit_20.fa_2  (    .a(\in_40<2> ),    .b(\in_41<2> ),    .cin(\adder_4bit_20.c<1> ),    .cout(\adder_4bit_20.c<2> ),    .s(\adder_4bit_20.s<2> )
  );
  full_adder \adder_4bit_20.fa_3  (    .a(\in_40<3> ),    .b(\in_41<3> ),    .cin(\adder_4bit_20.c<2> ),    .cout(\adder_4bit_20.c<3> ),    .s(\adder_4bit_20.s<3> )
  );
  adder_sign_extension \adder_4bit_20.fa_4  (    .a(\in_40<3> ),    .b(\in_41<3> ),    .cin(\adder_4bit_20.c<3> ),    .s(\adder_4bit_20.s<4> ),    .sign(sign_weight)
  );
  half_adder \adder_4bit_20.ha_0  (    .a(\in_40<0> ),    .b(\in_41<0> ),    .cout(\adder_4bit_20.c<0> ),    .s(\adder_4bit_20.s<0> )
  );
  full_adder \adder_4bit_21.fa_1  (    .a(\in_42<1> ),    .b(\in_43<1> ),    .cin(\adder_4bit_21.c<0> ),    .cout(\adder_4bit_21.c<1> ),    .s(\adder_4bit_21.s<1> )
  );
  full_adder \adder_4bit_21.fa_2  (    .a(\in_42<2> ),    .b(\in_43<2> ),    .cin(\adder_4bit_21.c<1> ),    .cout(\adder_4bit_21.c<2> ),    .s(\adder_4bit_21.s<2> )
  );
  full_adder \adder_4bit_21.fa_3  (    .a(\in_42<3> ),    .b(\in_43<3> ),    .cin(\adder_4bit_21.c<2> ),    .cout(\adder_4bit_21.c<3> ),    .s(\adder_4bit_21.s<3> )
  );
  adder_sign_extension \adder_4bit_21.fa_4  (    .a(\in_42<3> ),    .b(\in_43<3> ),    .cin(\adder_4bit_21.c<3> ),    .s(\adder_4bit_21.s<4> ),    .sign(sign_weight)
  );
  half_adder \adder_4bit_21.ha_0  (    .a(\in_42<0> ),    .b(\in_43<0> ),    .cout(\adder_4bit_21.c<0> ),    .s(\adder_4bit_21.s<0> )
  );
  full_adder \adder_4bit_22.fa_1  (    .a(\in_44<1> ),    .b(\in_45<1> ),    .cin(\adder_4bit_22.c<0> ),    .cout(\adder_4bit_22.c<1> ),    .s(\adder_4bit_22.s<1> )
  );
  full_adder \adder_4bit_22.fa_2  (    .a(\in_44<2> ),    .b(\in_45<2> ),    .cin(\adder_4bit_22.c<1> ),    .cout(\adder_4bit_22.c<2> ),    .s(\adder_4bit_22.s<2> )
  );
  full_adder \adder_4bit_22.fa_3  (    .a(\in_44<3> ),    .b(\in_45<3> ),    .cin(\adder_4bit_22.c<2> ),    .cout(\adder_4bit_22.c<3> ),    .s(\adder_4bit_22.s<3> )
  );
  adder_sign_extension \adder_4bit_22.fa_4  (    .a(\in_44<3> ),    .b(\in_45<3> ),    .cin(\adder_4bit_22.c<3> ),    .s(\adder_4bit_22.s<4> ),    .sign(sign_weight)
  );
  half_adder \adder_4bit_22.ha_0  (    .a(\in_44<0> ),    .b(\in_45<0> ),    .cout(\adder_4bit_22.c<0> ),    .s(\adder_4bit_22.s<0> )
  );
  full_adder \adder_4bit_23.fa_1  (    .a(\in_46<1> ),    .b(\in_47<1> ),    .cin(\adder_4bit_23.c<0> ),    .cout(\adder_4bit_23.c<1> ),    .s(\adder_4bit_23.s<1> )
  );
  full_adder \adder_4bit_23.fa_2  (    .a(\in_46<2> ),    .b(\in_47<2> ),    .cin(\adder_4bit_23.c<1> ),    .cout(\adder_4bit_23.c<2> ),    .s(\adder_4bit_23.s<2> )
  );
  full_adder \adder_4bit_23.fa_3  (    .a(\in_46<3> ),    .b(\in_47<3> ),    .cin(\adder_4bit_23.c<2> ),    .cout(\adder_4bit_23.c<3> ),    .s(\adder_4bit_23.s<3> )
  );
  adder_sign_extension \adder_4bit_23.fa_4  (    .a(\in_46<3> ),    .b(\in_47<3> ),    .cin(\adder_4bit_23.c<3> ),    .s(\adder_4bit_23.s<4> ),    .sign(sign_weight)
  );
  half_adder \adder_4bit_23.ha_0  (    .a(\in_46<0> ),    .b(\in_47<0> ),    .cout(\adder_4bit_23.c<0> ),    .s(\adder_4bit_23.s<0> )
  );
  full_adder \adder_4bit_24.fa_1  (    .a(\in_48<1> ),    .b(\in_49<1> ),    .cin(\adder_4bit_24.c<0> ),    .cout(\adder_4bit_24.c<1> ),    .s(\adder_4bit_24.s<1> )
  );
  full_adder \adder_4bit_24.fa_2  (    .a(\in_48<2> ),    .b(\in_49<2> ),    .cin(\adder_4bit_24.c<1> ),    .cout(\adder_4bit_24.c<2> ),    .s(\adder_4bit_24.s<2> )
  );
  full_adder \adder_4bit_24.fa_3  (    .a(\in_48<3> ),    .b(\in_49<3> ),    .cin(\adder_4bit_24.c<2> ),    .cout(\adder_4bit_24.c<3> ),    .s(\adder_4bit_24.s<3> )
  );
  adder_sign_extension \adder_4bit_24.fa_4  (    .a(\in_48<3> ),    .b(\in_49<3> ),    .cin(\adder_4bit_24.c<3> ),    .s(\adder_4bit_24.s<4> ),    .sign(sign_weight)
  );
  half_adder \adder_4bit_24.ha_0  (    .a(\in_48<0> ),    .b(\in_49<0> ),    .cout(\adder_4bit_24.c<0> ),    .s(\adder_4bit_24.s<0> )
  );
  full_adder \adder_4bit_25.fa_1  (    .a(\in_50<1> ),    .b(\in_51<1> ),    .cin(\adder_4bit_25.c<0> ),    .cout(\adder_4bit_25.c<1> ),    .s(\adder_4bit_25.s<1> )
  );
  full_adder \adder_4bit_25.fa_2  (    .a(\in_50<2> ),    .b(\in_51<2> ),    .cin(\adder_4bit_25.c<1> ),    .cout(\adder_4bit_25.c<2> ),    .s(\adder_4bit_25.s<2> )
  );
  full_adder \adder_4bit_25.fa_3  (    .a(\in_50<3> ),    .b(\in_51<3> ),    .cin(\adder_4bit_25.c<2> ),    .cout(\adder_4bit_25.c<3> ),    .s(\adder_4bit_25.s<3> )
  );
  adder_sign_extension \adder_4bit_25.fa_4  (    .a(\in_50<3> ),    .b(\in_51<3> ),    .cin(\adder_4bit_25.c<3> ),    .s(\adder_4bit_25.s<4> ),    .sign(sign_weight)
  );
  half_adder \adder_4bit_25.ha_0  (    .a(\in_50<0> ),    .b(\in_51<0> ),    .cout(\adder_4bit_25.c<0> ),    .s(\adder_4bit_25.s<0> )
  );
  full_adder \adder_4bit_26.fa_1  (    .a(\in_52<1> ),    .b(\in_53<1> ),    .cin(\adder_4bit_26.c<0> ),    .cout(\adder_4bit_26.c<1> ),    .s(\adder_4bit_26.s<1> )
  );
  full_adder \adder_4bit_26.fa_2  (    .a(\in_52<2> ),    .b(\in_53<2> ),    .cin(\adder_4bit_26.c<1> ),    .cout(\adder_4bit_26.c<2> ),    .s(\adder_4bit_26.s<2> )
  );
  full_adder \adder_4bit_26.fa_3  (    .a(\in_52<3> ),    .b(\in_53<3> ),    .cin(\adder_4bit_26.c<2> ),    .cout(\adder_4bit_26.c<3> ),    .s(\adder_4bit_26.s<3> )
  );
  adder_sign_extension \adder_4bit_26.fa_4  (    .a(\in_52<3> ),    .b(\in_53<3> ),    .cin(\adder_4bit_26.c<3> ),    .s(\adder_4bit_26.s<4> ),    .sign(sign_weight)
  );
  half_adder \adder_4bit_26.ha_0  (    .a(\in_52<0> ),    .b(\in_53<0> ),    .cout(\adder_4bit_26.c<0> ),    .s(\adder_4bit_26.s<0> )
  );
  full_adder \adder_4bit_27.fa_1  (    .a(\in_54<1> ),    .b(\in_55<1> ),    .cin(\adder_4bit_27.c<0> ),    .cout(\adder_4bit_27.c<1> ),    .s(\adder_4bit_27.s<1> )
  );
  full_adder \adder_4bit_27.fa_2  (    .a(\in_54<2> ),    .b(\in_55<2> ),    .cin(\adder_4bit_27.c<1> ),    .cout(\adder_4bit_27.c<2> ),    .s(\adder_4bit_27.s<2> )
  );
  full_adder \adder_4bit_27.fa_3  (    .a(\in_54<3> ),    .b(\in_55<3> ),    .cin(\adder_4bit_27.c<2> ),    .cout(\adder_4bit_27.c<3> ),    .s(\adder_4bit_27.s<3> )
  );
  adder_sign_extension \adder_4bit_27.fa_4  (    .a(\in_54<3> ),    .b(\in_55<3> ),    .cin(\adder_4bit_27.c<3> ),    .s(\adder_4bit_27.s<4> ),    .sign(sign_weight)
  );
  half_adder \adder_4bit_27.ha_0  (    .a(\in_54<0> ),    .b(\in_55<0> ),    .cout(\adder_4bit_27.c<0> ),    .s(\adder_4bit_27.s<0> )
  );
  full_adder \adder_4bit_28.fa_1  (    .a(\in_56<1> ),    .b(\in_57<1> ),    .cin(\adder_4bit_28.c<0> ),    .cout(\adder_4bit_28.c<1> ),    .s(\adder_4bit_28.s<1> )
  );
  full_adder \adder_4bit_28.fa_2  (    .a(\in_56<2> ),    .b(\in_57<2> ),    .cin(\adder_4bit_28.c<1> ),    .cout(\adder_4bit_28.c<2> ),    .s(\adder_4bit_28.s<2> )
  );
  full_adder \adder_4bit_28.fa_3  (    .a(\in_56<3> ),    .b(\in_57<3> ),    .cin(\adder_4bit_28.c<2> ),    .cout(\adder_4bit_28.c<3> ),    .s(\adder_4bit_28.s<3> )
  );
  adder_sign_extension \adder_4bit_28.fa_4  (    .a(\in_56<3> ),    .b(\in_57<3> ),    .cin(\adder_4bit_28.c<3> ),    .s(\adder_4bit_28.s<4> ),    .sign(sign_weight)
  );
  half_adder \adder_4bit_28.ha_0  (    .a(\in_56<0> ),    .b(\in_57<0> ),    .cout(\adder_4bit_28.c<0> ),    .s(\adder_4bit_28.s<0> )
  );
  full_adder \adder_4bit_29.fa_1  (    .a(\in_58<1> ),    .b(\in_59<1> ),    .cin(\adder_4bit_29.c<0> ),    .cout(\adder_4bit_29.c<1> ),    .s(\adder_4bit_29.s<1> )
  );
  full_adder \adder_4bit_29.fa_2  (    .a(\in_58<2> ),    .b(\in_59<2> ),    .cin(\adder_4bit_29.c<1> ),    .cout(\adder_4bit_29.c<2> ),    .s(\adder_4bit_29.s<2> )
  );
  full_adder \adder_4bit_29.fa_3  (    .a(\in_58<3> ),    .b(\in_59<3> ),    .cin(\adder_4bit_29.c<2> ),    .cout(\adder_4bit_29.c<3> ),    .s(\adder_4bit_29.s<3> )
  );
  adder_sign_extension \adder_4bit_29.fa_4  (    .a(\in_58<3> ),    .b(\in_59<3> ),    .cin(\adder_4bit_29.c<3> ),    .s(\adder_4bit_29.s<4> ),    .sign(sign_weight)
  );
  half_adder \adder_4bit_29.ha_0  (    .a(\in_58<0> ),    .b(\in_59<0> ),    .cout(\adder_4bit_29.c<0> ),    .s(\adder_4bit_29.s<0> )
  );
  full_adder \adder_4bit_3.fa_1  (    .a(\in_6<1> ),    .b(\in_7<1> ),    .cin(\adder_4bit_3.c<0> ),    .cout(\adder_4bit_3.c<1> ),    .s(\adder_4bit_3.s<1> )
  );
  full_adder \adder_4bit_3.fa_2  (    .a(\in_6<2> ),    .b(\in_7<2> ),    .cin(\adder_4bit_3.c<1> ),    .cout(\adder_4bit_3.c<2> ),    .s(\adder_4bit_3.s<2> )
  );
  full_adder \adder_4bit_3.fa_3  (    .a(\in_6<3> ),    .b(\in_7<3> ),    .cin(\adder_4bit_3.c<2> ),    .cout(\adder_4bit_3.c<3> ),    .s(\adder_4bit_3.s<3> )
  );
  adder_sign_extension \adder_4bit_3.fa_4  (    .a(\in_6<3> ),    .b(\in_7<3> ),    .cin(\adder_4bit_3.c<3> ),    .s(\adder_4bit_3.s<4> ),    .sign(sign_weight)
  );
  half_adder \adder_4bit_3.ha_0  (    .a(\in_6<0> ),    .b(\in_7<0> ),    .cout(\adder_4bit_3.c<0> ),    .s(\adder_4bit_3.s<0> )
  );
  full_adder \adder_4bit_30.fa_1  (    .a(\in_60<1> ),    .b(\in_61<1> ),    .cin(\adder_4bit_30.c<0> ),    .cout(\adder_4bit_30.c<1> ),    .s(\adder_4bit_30.s<1> )
  );
  full_adder \adder_4bit_30.fa_2  (    .a(\in_60<2> ),    .b(\in_61<2> ),    .cin(\adder_4bit_30.c<1> ),    .cout(\adder_4bit_30.c<2> ),    .s(\adder_4bit_30.s<2> )
  );
  full_adder \adder_4bit_30.fa_3  (    .a(\in_60<3> ),    .b(\in_61<3> ),    .cin(\adder_4bit_30.c<2> ),    .cout(\adder_4bit_30.c<3> ),    .s(\adder_4bit_30.s<3> )
  );
  adder_sign_extension \adder_4bit_30.fa_4  (    .a(\in_60<3> ),    .b(\in_61<3> ),    .cin(\adder_4bit_30.c<3> ),    .s(\adder_4bit_30.s<4> ),    .sign(sign_weight)
  );
  half_adder \adder_4bit_30.ha_0  (    .a(\in_60<0> ),    .b(\in_61<0> ),    .cout(\adder_4bit_30.c<0> ),    .s(\adder_4bit_30.s<0> )
  );
  full_adder \adder_4bit_31.fa_1  (    .a(\in_62<1> ),    .b(\in_63<1> ),    .cin(\adder_4bit_31.c<0> ),    .cout(\adder_4bit_31.c<1> ),    .s(\adder_4bit_31.s<1> )
  );
  full_adder \adder_4bit_31.fa_2  (    .a(\in_62<2> ),    .b(\in_63<2> ),    .cin(\adder_4bit_31.c<1> ),    .cout(\adder_4bit_31.c<2> ),    .s(\adder_4bit_31.s<2> )
  );
  full_adder \adder_4bit_31.fa_3  (    .a(\in_62<3> ),    .b(\in_63<3> ),    .cin(\adder_4bit_31.c<2> ),    .cout(\adder_4bit_31.c<3> ),    .s(\adder_4bit_31.s<3> )
  );
  adder_sign_extension \adder_4bit_31.fa_4  (    .a(\in_62<3> ),    .b(\in_63<3> ),    .cin(\adder_4bit_31.c<3> ),    .s(\adder_4bit_31.s<4> ),    .sign(sign_weight)
  );
  half_adder \adder_4bit_31.ha_0  (    .a(\in_62<0> ),    .b(\in_63<0> ),    .cout(\adder_4bit_31.c<0> ),    .s(\adder_4bit_31.s<0> )
  );
  full_adder \adder_4bit_4.fa_1  (    .a(\in_8<1> ),    .b(\in_9<1> ),    .cin(\adder_4bit_4.c<0> ),    .cout(\adder_4bit_4.c<1> ),    .s(\adder_4bit_4.s<1> )
  );
  full_adder \adder_4bit_4.fa_2  (    .a(\in_8<2> ),    .b(\in_9<2> ),    .cin(\adder_4bit_4.c<1> ),    .cout(\adder_4bit_4.c<2> ),    .s(\adder_4bit_4.s<2> )
  );
  full_adder \adder_4bit_4.fa_3  (    .a(\in_8<3> ),    .b(\in_9<3> ),    .cin(\adder_4bit_4.c<2> ),    .cout(\adder_4bit_4.c<3> ),    .s(\adder_4bit_4.s<3> )
  );
  adder_sign_extension \adder_4bit_4.fa_4  (    .a(\in_8<3> ),    .b(\in_9<3> ),    .cin(\adder_4bit_4.c<3> ),    .s(\adder_4bit_4.s<4> ),    .sign(sign_weight)
  );
  half_adder \adder_4bit_4.ha_0  (    .a(\in_8<0> ),    .b(\in_9<0> ),    .cout(\adder_4bit_4.c<0> ),    .s(\adder_4bit_4.s<0> )
  );
  full_adder \adder_4bit_5.fa_1  (    .a(\in_10<1> ),    .b(\in_11<1> ),    .cin(\adder_4bit_5.c<0> ),    .cout(\adder_4bit_5.c<1> ),    .s(\adder_4bit_5.s<1> )
  );
  full_adder \adder_4bit_5.fa_2  (    .a(\in_10<2> ),    .b(\in_11<2> ),    .cin(\adder_4bit_5.c<1> ),    .cout(\adder_4bit_5.c<2> ),    .s(\adder_4bit_5.s<2> )
  );
  full_adder \adder_4bit_5.fa_3  (    .a(\in_10<3> ),    .b(\in_11<3> ),    .cin(\adder_4bit_5.c<2> ),    .cout(\adder_4bit_5.c<3> ),    .s(\adder_4bit_5.s<3> )
  );
  adder_sign_extension \adder_4bit_5.fa_4  (    .a(\in_10<3> ),    .b(\in_11<3> ),    .cin(\adder_4bit_5.c<3> ),    .s(\adder_4bit_5.s<4> ),    .sign(sign_weight)
  );
  half_adder \adder_4bit_5.ha_0  (    .a(\in_10<0> ),    .b(\in_11<0> ),    .cout(\adder_4bit_5.c<0> ),    .s(\adder_4bit_5.s<0> )
  );
  full_adder \adder_4bit_6.fa_1  (    .a(\in_12<1> ),    .b(\in_13<1> ),    .cin(\adder_4bit_6.c<0> ),    .cout(\adder_4bit_6.c<1> ),    .s(\adder_4bit_6.s<1> )
  );
  full_adder \adder_4bit_6.fa_2  (    .a(\in_12<2> ),    .b(\in_13<2> ),    .cin(\adder_4bit_6.c<1> ),    .cout(\adder_4bit_6.c<2> ),    .s(\adder_4bit_6.s<2> )
  );
  full_adder \adder_4bit_6.fa_3  (    .a(\in_12<3> ),    .b(\in_13<3> ),    .cin(\adder_4bit_6.c<2> ),    .cout(\adder_4bit_6.c<3> ),    .s(\adder_4bit_6.s<3> )
  );
  adder_sign_extension \adder_4bit_6.fa_4  (    .a(\in_12<3> ),    .b(\in_13<3> ),    .cin(\adder_4bit_6.c<3> ),    .s(\adder_4bit_6.s<4> ),    .sign(sign_weight)
  );
  half_adder \adder_4bit_6.ha_0  (    .a(\in_12<0> ),    .b(\in_13<0> ),    .cout(\adder_4bit_6.c<0> ),    .s(\adder_4bit_6.s<0> )
  );
  full_adder \adder_4bit_7.fa_1  (    .a(\in_14<1> ),    .b(\in_15<1> ),    .cin(\adder_4bit_7.c<0> ),    .cout(\adder_4bit_7.c<1> ),    .s(\adder_4bit_7.s<1> )
  );
  full_adder \adder_4bit_7.fa_2  (    .a(\in_14<2> ),    .b(\in_15<2> ),    .cin(\adder_4bit_7.c<1> ),    .cout(\adder_4bit_7.c<2> ),    .s(\adder_4bit_7.s<2> )
  );
  full_adder \adder_4bit_7.fa_3  (    .a(\in_14<3> ),    .b(\in_15<3> ),    .cin(\adder_4bit_7.c<2> ),    .cout(\adder_4bit_7.c<3> ),    .s(\adder_4bit_7.s<3> )
  );
  adder_sign_extension \adder_4bit_7.fa_4  (    .a(\in_14<3> ),    .b(\in_15<3> ),    .cin(\adder_4bit_7.c<3> ),    .s(\adder_4bit_7.s<4> ),    .sign(sign_weight)
  );
  half_adder \adder_4bit_7.ha_0  (    .a(\in_14<0> ),    .b(\in_15<0> ),    .cout(\adder_4bit_7.c<0> ),    .s(\adder_4bit_7.s<0> )
  );
  full_adder \adder_4bit_8.fa_1  (    .a(\in_16<1> ),    .b(\in_17<1> ),    .cin(\adder_4bit_8.c<0> ),    .cout(\adder_4bit_8.c<1> ),    .s(\adder_4bit_8.s<1> )
  );
  full_adder \adder_4bit_8.fa_2  (    .a(\in_16<2> ),    .b(\in_17<2> ),    .cin(\adder_4bit_8.c<1> ),    .cout(\adder_4bit_8.c<2> ),    .s(\adder_4bit_8.s<2> )
  );
  full_adder \adder_4bit_8.fa_3  (    .a(\in_16<3> ),    .b(\in_17<3> ),    .cin(\adder_4bit_8.c<2> ),    .cout(\adder_4bit_8.c<3> ),    .s(\adder_4bit_8.s<3> )
  );
  adder_sign_extension \adder_4bit_8.fa_4  (    .a(\in_16<3> ),    .b(\in_17<3> ),    .cin(\adder_4bit_8.c<3> ),    .s(\adder_4bit_8.s<4> ),    .sign(sign_weight)
  );
  half_adder \adder_4bit_8.ha_0  (    .a(\in_16<0> ),    .b(\in_17<0> ),    .cout(\adder_4bit_8.c<0> ),    .s(\adder_4bit_8.s<0> )
  );
  full_adder \adder_4bit_9.fa_1  (    .a(\in_18<1> ),    .b(\in_19<1> ),    .cin(\adder_4bit_9.c<0> ),    .cout(\adder_4bit_9.c<1> ),    .s(\adder_4bit_9.s<1> )
  );
  full_adder \adder_4bit_9.fa_2  (    .a(\in_18<2> ),    .b(\in_19<2> ),    .cin(\adder_4bit_9.c<1> ),    .cout(\adder_4bit_9.c<2> ),    .s(\adder_4bit_9.s<2> )
  );
  full_adder \adder_4bit_9.fa_3  (    .a(\in_18<3> ),    .b(\in_19<3> ),    .cin(\adder_4bit_9.c<2> ),    .cout(\adder_4bit_9.c<3> ),    .s(\adder_4bit_9.s<3> )
  );
  adder_sign_extension \adder_4bit_9.fa_4  (    .a(\in_18<3> ),    .b(\in_19<3> ),    .cin(\adder_4bit_9.c<3> ),    .s(\adder_4bit_9.s<4> ),    .sign(sign_weight)
  );
  half_adder \adder_4bit_9.ha_0  (    .a(\in_18<0> ),    .b(\in_19<0> ),    .cout(\adder_4bit_9.c<0> ),    .s(\adder_4bit_9.s<0> )
  );
  full_adder \adder_5bit_0.fa_1  (    .a(\adder_4bit_0.s<1> ),    .b(\adder_4bit_1.s<1> ),    .cin(\adder_5bit_0.c<0> ),    .cout(\adder_5bit_0.c<1> ),    .s(\adder_5bit_0.s<1> )
  );
  full_adder \adder_5bit_0.fa_2  (    .a(\adder_4bit_0.s<2> ),    .b(\adder_4bit_1.s<2> ),    .cin(\adder_5bit_0.c<1> ),    .cout(\adder_5bit_0.c<2> ),    .s(\adder_5bit_0.s<2> )
  );
  full_adder \adder_5bit_0.fa_3  (    .a(\adder_4bit_0.s<3> ),    .b(\adder_4bit_1.s<3> ),    .cin(\adder_5bit_0.c<2> ),    .cout(\adder_5bit_0.c<3> ),    .s(\adder_5bit_0.s<3> )
  );
  full_adder \adder_5bit_0.fa_4  (    .a(\adder_4bit_0.s<4> ),    .b(\adder_4bit_1.s<4> ),    .cin(\adder_5bit_0.c<3> ),    .cout(\adder_5bit_0.c<4> ),    .s(\adder_5bit_0.s<4> )
  );
  adder_sign_extension \adder_5bit_0.fa_5  (    .a(\adder_4bit_0.s<4> ),    .b(\adder_4bit_1.s<4> ),    .cin(\adder_5bit_0.c<4> ),    .s(\adder_5bit_0.s<5> ),    .sign(sign_weight)
  );
  half_adder \adder_5bit_0.ha_0  (    .a(\adder_4bit_0.s<0> ),    .b(\adder_4bit_1.s<0> ),    .cout(\adder_5bit_0.c<0> ),    .s(\adder_5bit_0.s<0> )
  );
  full_adder \adder_5bit_1.fa_1  (    .a(\adder_4bit_2.s<1> ),    .b(\adder_4bit_3.s<1> ),    .cin(\adder_5bit_1.c<0> ),    .cout(\adder_5bit_1.c<1> ),    .s(\adder_5bit_1.s<1> )
  );
  full_adder \adder_5bit_1.fa_2  (    .a(\adder_4bit_2.s<2> ),    .b(\adder_4bit_3.s<2> ),    .cin(\adder_5bit_1.c<1> ),    .cout(\adder_5bit_1.c<2> ),    .s(\adder_5bit_1.s<2> )
  );
  full_adder \adder_5bit_1.fa_3  (    .a(\adder_4bit_2.s<3> ),    .b(\adder_4bit_3.s<3> ),    .cin(\adder_5bit_1.c<2> ),    .cout(\adder_5bit_1.c<3> ),    .s(\adder_5bit_1.s<3> )
  );
  full_adder \adder_5bit_1.fa_4  (    .a(\adder_4bit_2.s<4> ),    .b(\adder_4bit_3.s<4> ),    .cin(\adder_5bit_1.c<3> ),    .cout(\adder_5bit_1.c<4> ),    .s(\adder_5bit_1.s<4> )
  );
  adder_sign_extension \adder_5bit_1.fa_5  (    .a(\adder_4bit_2.s<4> ),    .b(\adder_4bit_3.s<4> ),    .cin(\adder_5bit_1.c<4> ),    .s(\adder_5bit_1.s<5> ),    .sign(sign_weight)
  );
  half_adder \adder_5bit_1.ha_0  (    .a(\adder_4bit_2.s<0> ),    .b(\adder_4bit_3.s<0> ),    .cout(\adder_5bit_1.c<0> ),    .s(\adder_5bit_1.s<0> )
  );
  full_adder \adder_5bit_10.fa_1  (    .a(\adder_4bit_20.s<1> ),    .b(\adder_4bit_21.s<1> ),    .cin(\adder_5bit_10.c<0> ),    .cout(\adder_5bit_10.c<1> ),    .s(\adder_5bit_10.s<1> )
  );
  full_adder \adder_5bit_10.fa_2  (    .a(\adder_4bit_20.s<2> ),    .b(\adder_4bit_21.s<2> ),    .cin(\adder_5bit_10.c<1> ),    .cout(\adder_5bit_10.c<2> ),    .s(\adder_5bit_10.s<2> )
  );
  full_adder \adder_5bit_10.fa_3  (    .a(\adder_4bit_20.s<3> ),    .b(\adder_4bit_21.s<3> ),    .cin(\adder_5bit_10.c<2> ),    .cout(\adder_5bit_10.c<3> ),    .s(\adder_5bit_10.s<3> )
  );
  full_adder \adder_5bit_10.fa_4  (    .a(\adder_4bit_20.s<4> ),    .b(\adder_4bit_21.s<4> ),    .cin(\adder_5bit_10.c<3> ),    .cout(\adder_5bit_10.c<4> ),    .s(\adder_5bit_10.s<4> )
  );
  adder_sign_extension \adder_5bit_10.fa_5  (    .a(\adder_4bit_20.s<4> ),    .b(\adder_4bit_21.s<4> ),    .cin(\adder_5bit_10.c<4> ),    .s(\adder_5bit_10.s<5> ),    .sign(sign_weight)
  );
  half_adder \adder_5bit_10.ha_0  (    .a(\adder_4bit_20.s<0> ),    .b(\adder_4bit_21.s<0> ),    .cout(\adder_5bit_10.c<0> ),    .s(\adder_5bit_10.s<0> )
  );
  full_adder \adder_5bit_11.fa_1  (    .a(\adder_4bit_22.s<1> ),    .b(\adder_4bit_23.s<1> ),    .cin(\adder_5bit_11.c<0> ),    .cout(\adder_5bit_11.c<1> ),    .s(\adder_5bit_11.s<1> )
  );
  full_adder \adder_5bit_11.fa_2  (    .a(\adder_4bit_22.s<2> ),    .b(\adder_4bit_23.s<2> ),    .cin(\adder_5bit_11.c<1> ),    .cout(\adder_5bit_11.c<2> ),    .s(\adder_5bit_11.s<2> )
  );
  full_adder \adder_5bit_11.fa_3  (    .a(\adder_4bit_22.s<3> ),    .b(\adder_4bit_23.s<3> ),    .cin(\adder_5bit_11.c<2> ),    .cout(\adder_5bit_11.c<3> ),    .s(\adder_5bit_11.s<3> )
  );
  full_adder \adder_5bit_11.fa_4  (    .a(\adder_4bit_22.s<4> ),    .b(\adder_4bit_23.s<4> ),    .cin(\adder_5bit_11.c<3> ),    .cout(\adder_5bit_11.c<4> ),    .s(\adder_5bit_11.s<4> )
  );
  adder_sign_extension \adder_5bit_11.fa_5  (    .a(\adder_4bit_22.s<4> ),    .b(\adder_4bit_23.s<4> ),    .cin(\adder_5bit_11.c<4> ),    .s(\adder_5bit_11.s<5> ),    .sign(sign_weight)
  );
  half_adder \adder_5bit_11.ha_0  (    .a(\adder_4bit_22.s<0> ),    .b(\adder_4bit_23.s<0> ),    .cout(\adder_5bit_11.c<0> ),    .s(\adder_5bit_11.s<0> )
  );
  full_adder \adder_5bit_12.fa_1  (    .a(\adder_4bit_24.s<1> ),    .b(\adder_4bit_25.s<1> ),    .cin(\adder_5bit_12.c<0> ),    .cout(\adder_5bit_12.c<1> ),    .s(\adder_5bit_12.s<1> )
  );
  full_adder \adder_5bit_12.fa_2  (    .a(\adder_4bit_24.s<2> ),    .b(\adder_4bit_25.s<2> ),    .cin(\adder_5bit_12.c<1> ),    .cout(\adder_5bit_12.c<2> ),    .s(\adder_5bit_12.s<2> )
  );
  full_adder \adder_5bit_12.fa_3  (    .a(\adder_4bit_24.s<3> ),    .b(\adder_4bit_25.s<3> ),    .cin(\adder_5bit_12.c<2> ),    .cout(\adder_5bit_12.c<3> ),    .s(\adder_5bit_12.s<3> )
  );
  full_adder \adder_5bit_12.fa_4  (    .a(\adder_4bit_24.s<4> ),    .b(\adder_4bit_25.s<4> ),    .cin(\adder_5bit_12.c<3> ),    .cout(\adder_5bit_12.c<4> ),    .s(\adder_5bit_12.s<4> )
  );
  adder_sign_extension \adder_5bit_12.fa_5  (    .a(\adder_4bit_24.s<4> ),    .b(\adder_4bit_25.s<4> ),    .cin(\adder_5bit_12.c<4> ),    .s(\adder_5bit_12.s<5> ),    .sign(sign_weight)
  );
  half_adder \adder_5bit_12.ha_0  (    .a(\adder_4bit_24.s<0> ),    .b(\adder_4bit_25.s<0> ),    .cout(\adder_5bit_12.c<0> ),    .s(\adder_5bit_12.s<0> )
  );
  full_adder \adder_5bit_13.fa_1  (    .a(\adder_4bit_26.s<1> ),    .b(\adder_4bit_27.s<1> ),    .cin(\adder_5bit_13.c<0> ),    .cout(\adder_5bit_13.c<1> ),    .s(\adder_5bit_13.s<1> )
  );
  full_adder \adder_5bit_13.fa_2  (    .a(\adder_4bit_26.s<2> ),    .b(\adder_4bit_27.s<2> ),    .cin(\adder_5bit_13.c<1> ),    .cout(\adder_5bit_13.c<2> ),    .s(\adder_5bit_13.s<2> )
  );
  full_adder \adder_5bit_13.fa_3  (    .a(\adder_4bit_26.s<3> ),    .b(\adder_4bit_27.s<3> ),    .cin(\adder_5bit_13.c<2> ),    .cout(\adder_5bit_13.c<3> ),    .s(\adder_5bit_13.s<3> )
  );
  full_adder \adder_5bit_13.fa_4  (    .a(\adder_4bit_26.s<4> ),    .b(\adder_4bit_27.s<4> ),    .cin(\adder_5bit_13.c<3> ),    .cout(\adder_5bit_13.c<4> ),    .s(\adder_5bit_13.s<4> )
  );
  adder_sign_extension \adder_5bit_13.fa_5  (    .a(\adder_4bit_26.s<4> ),    .b(\adder_4bit_27.s<4> ),    .cin(\adder_5bit_13.c<4> ),    .s(\adder_5bit_13.s<5> ),    .sign(sign_weight)
  );
  half_adder \adder_5bit_13.ha_0  (    .a(\adder_4bit_26.s<0> ),    .b(\adder_4bit_27.s<0> ),    .cout(\adder_5bit_13.c<0> ),    .s(\adder_5bit_13.s<0> )
  );
  full_adder \adder_5bit_14.fa_1  (    .a(\adder_4bit_28.s<1> ),    .b(\adder_4bit_29.s<1> ),    .cin(\adder_5bit_14.c<0> ),    .cout(\adder_5bit_14.c<1> ),    .s(\adder_5bit_14.s<1> )
  );
  full_adder \adder_5bit_14.fa_2  (    .a(\adder_4bit_28.s<2> ),    .b(\adder_4bit_29.s<2> ),    .cin(\adder_5bit_14.c<1> ),    .cout(\adder_5bit_14.c<2> ),    .s(\adder_5bit_14.s<2> )
  );
  full_adder \adder_5bit_14.fa_3  (    .a(\adder_4bit_28.s<3> ),    .b(\adder_4bit_29.s<3> ),    .cin(\adder_5bit_14.c<2> ),    .cout(\adder_5bit_14.c<3> ),    .s(\adder_5bit_14.s<3> )
  );
  full_adder \adder_5bit_14.fa_4  (    .a(\adder_4bit_28.s<4> ),    .b(\adder_4bit_29.s<4> ),    .cin(\adder_5bit_14.c<3> ),    .cout(\adder_5bit_14.c<4> ),    .s(\adder_5bit_14.s<4> )
  );
  adder_sign_extension \adder_5bit_14.fa_5  (    .a(\adder_4bit_28.s<4> ),    .b(\adder_4bit_29.s<4> ),    .cin(\adder_5bit_14.c<4> ),    .s(\adder_5bit_14.s<5> ),    .sign(sign_weight)
  );
  half_adder \adder_5bit_14.ha_0  (    .a(\adder_4bit_28.s<0> ),    .b(\adder_4bit_29.s<0> ),    .cout(\adder_5bit_14.c<0> ),    .s(\adder_5bit_14.s<0> )
  );
  full_adder \adder_5bit_15.fa_1  (    .a(\adder_4bit_30.s<1> ),    .b(\adder_4bit_31.s<1> ),    .cin(\adder_5bit_15.c<0> ),    .cout(\adder_5bit_15.c<1> ),    .s(\adder_5bit_15.s<1> )
  );
  full_adder \adder_5bit_15.fa_2  (    .a(\adder_4bit_30.s<2> ),    .b(\adder_4bit_31.s<2> ),    .cin(\adder_5bit_15.c<1> ),    .cout(\adder_5bit_15.c<2> ),    .s(\adder_5bit_15.s<2> )
  );
  full_adder \adder_5bit_15.fa_3  (    .a(\adder_4bit_30.s<3> ),    .b(\adder_4bit_31.s<3> ),    .cin(\adder_5bit_15.c<2> ),    .cout(\adder_5bit_15.c<3> ),    .s(\adder_5bit_15.s<3> )
  );
  full_adder \adder_5bit_15.fa_4  (    .a(\adder_4bit_30.s<4> ),    .b(\adder_4bit_31.s<4> ),    .cin(\adder_5bit_15.c<3> ),    .cout(\adder_5bit_15.c<4> ),    .s(\adder_5bit_15.s<4> )
  );
  adder_sign_extension \adder_5bit_15.fa_5  (    .a(\adder_4bit_30.s<4> ),    .b(\adder_4bit_31.s<4> ),    .cin(\adder_5bit_15.c<4> ),    .s(\adder_5bit_15.s<5> ),    .sign(sign_weight)
  );
  half_adder \adder_5bit_15.ha_0  (    .a(\adder_4bit_30.s<0> ),    .b(\adder_4bit_31.s<0> ),    .cout(\adder_5bit_15.c<0> ),    .s(\adder_5bit_15.s<0> )
  );
  full_adder \adder_5bit_2.fa_1  (    .a(\adder_4bit_4.s<1> ),    .b(\adder_4bit_5.s<1> ),    .cin(\adder_5bit_2.c<0> ),    .cout(\adder_5bit_2.c<1> ),    .s(\adder_5bit_2.s<1> )
  );
  full_adder \adder_5bit_2.fa_2  (    .a(\adder_4bit_4.s<2> ),    .b(\adder_4bit_5.s<2> ),    .cin(\adder_5bit_2.c<1> ),    .cout(\adder_5bit_2.c<2> ),    .s(\adder_5bit_2.s<2> )
  );
  full_adder \adder_5bit_2.fa_3  (    .a(\adder_4bit_4.s<3> ),    .b(\adder_4bit_5.s<3> ),    .cin(\adder_5bit_2.c<2> ),    .cout(\adder_5bit_2.c<3> ),    .s(\adder_5bit_2.s<3> )
  );
  full_adder \adder_5bit_2.fa_4  (    .a(\adder_4bit_4.s<4> ),    .b(\adder_4bit_5.s<4> ),    .cin(\adder_5bit_2.c<3> ),    .cout(\adder_5bit_2.c<4> ),    .s(\adder_5bit_2.s<4> )
  );
  adder_sign_extension \adder_5bit_2.fa_5  (    .a(\adder_4bit_4.s<4> ),    .b(\adder_4bit_5.s<4> ),    .cin(\adder_5bit_2.c<4> ),    .s(\adder_5bit_2.s<5> ),    .sign(sign_weight)
  );
  half_adder \adder_5bit_2.ha_0  (    .a(\adder_4bit_4.s<0> ),    .b(\adder_4bit_5.s<0> ),    .cout(\adder_5bit_2.c<0> ),    .s(\adder_5bit_2.s<0> )
  );
  full_adder \adder_5bit_3.fa_1  (    .a(\adder_4bit_6.s<1> ),    .b(\adder_4bit_7.s<1> ),    .cin(\adder_5bit_3.c<0> ),    .cout(\adder_5bit_3.c<1> ),    .s(\adder_5bit_3.s<1> )
  );
  full_adder \adder_5bit_3.fa_2  (    .a(\adder_4bit_6.s<2> ),    .b(\adder_4bit_7.s<2> ),    .cin(\adder_5bit_3.c<1> ),    .cout(\adder_5bit_3.c<2> ),    .s(\adder_5bit_3.s<2> )
  );
  full_adder \adder_5bit_3.fa_3  (    .a(\adder_4bit_6.s<3> ),    .b(\adder_4bit_7.s<3> ),    .cin(\adder_5bit_3.c<2> ),    .cout(\adder_5bit_3.c<3> ),    .s(\adder_5bit_3.s<3> )
  );
  full_adder \adder_5bit_3.fa_4  (    .a(\adder_4bit_6.s<4> ),    .b(\adder_4bit_7.s<4> ),    .cin(\adder_5bit_3.c<3> ),    .cout(\adder_5bit_3.c<4> ),    .s(\adder_5bit_3.s<4> )
  );
  adder_sign_extension \adder_5bit_3.fa_5  (    .a(\adder_4bit_6.s<4> ),    .b(\adder_4bit_7.s<4> ),    .cin(\adder_5bit_3.c<4> ),    .s(\adder_5bit_3.s<5> ),    .sign(sign_weight)
  );
  half_adder \adder_5bit_3.ha_0  (    .a(\adder_4bit_6.s<0> ),    .b(\adder_4bit_7.s<0> ),    .cout(\adder_5bit_3.c<0> ),    .s(\adder_5bit_3.s<0> )
  );
  full_adder \adder_5bit_4.fa_1  (    .a(\adder_4bit_8.s<1> ),    .b(\adder_4bit_9.s<1> ),    .cin(\adder_5bit_4.c<0> ),    .cout(\adder_5bit_4.c<1> ),    .s(\adder_5bit_4.s<1> )
  );
  full_adder \adder_5bit_4.fa_2  (    .a(\adder_4bit_8.s<2> ),    .b(\adder_4bit_9.s<2> ),    .cin(\adder_5bit_4.c<1> ),    .cout(\adder_5bit_4.c<2> ),    .s(\adder_5bit_4.s<2> )
  );
  full_adder \adder_5bit_4.fa_3  (    .a(\adder_4bit_8.s<3> ),    .b(\adder_4bit_9.s<3> ),    .cin(\adder_5bit_4.c<2> ),    .cout(\adder_5bit_4.c<3> ),    .s(\adder_5bit_4.s<3> )
  );
  full_adder \adder_5bit_4.fa_4  (    .a(\adder_4bit_8.s<4> ),    .b(\adder_4bit_9.s<4> ),    .cin(\adder_5bit_4.c<3> ),    .cout(\adder_5bit_4.c<4> ),    .s(\adder_5bit_4.s<4> )
  );
  adder_sign_extension \adder_5bit_4.fa_5  (    .a(\adder_4bit_8.s<4> ),    .b(\adder_4bit_9.s<4> ),    .cin(\adder_5bit_4.c<4> ),    .s(\adder_5bit_4.s<5> ),    .sign(sign_weight)
  );
  half_adder \adder_5bit_4.ha_0  (    .a(\adder_4bit_8.s<0> ),    .b(\adder_4bit_9.s<0> ),    .cout(\adder_5bit_4.c<0> ),    .s(\adder_5bit_4.s<0> )
  );
  full_adder \adder_5bit_5.fa_1  (    .a(\adder_4bit_10.s<1> ),    .b(\adder_4bit_11.s<1> ),    .cin(\adder_5bit_5.c<0> ),    .cout(\adder_5bit_5.c<1> ),    .s(\adder_5bit_5.s<1> )
  );
  full_adder \adder_5bit_5.fa_2  (    .a(\adder_4bit_10.s<2> ),    .b(\adder_4bit_11.s<2> ),    .cin(\adder_5bit_5.c<1> ),    .cout(\adder_5bit_5.c<2> ),    .s(\adder_5bit_5.s<2> )
  );
  full_adder \adder_5bit_5.fa_3  (    .a(\adder_4bit_10.s<3> ),    .b(\adder_4bit_11.s<3> ),    .cin(\adder_5bit_5.c<2> ),    .cout(\adder_5bit_5.c<3> ),    .s(\adder_5bit_5.s<3> )
  );
  full_adder \adder_5bit_5.fa_4  (    .a(\adder_4bit_10.s<4> ),    .b(\adder_4bit_11.s<4> ),    .cin(\adder_5bit_5.c<3> ),    .cout(\adder_5bit_5.c<4> ),    .s(\adder_5bit_5.s<4> )
  );
  adder_sign_extension \adder_5bit_5.fa_5  (    .a(\adder_4bit_10.s<4> ),    .b(\adder_4bit_11.s<4> ),    .cin(\adder_5bit_5.c<4> ),    .s(\adder_5bit_5.s<5> ),    .sign(sign_weight)
  );
  half_adder \adder_5bit_5.ha_0  (    .a(\adder_4bit_10.s<0> ),    .b(\adder_4bit_11.s<0> ),    .cout(\adder_5bit_5.c<0> ),    .s(\adder_5bit_5.s<0> )
  );
  full_adder \adder_5bit_6.fa_1  (    .a(\adder_4bit_12.s<1> ),    .b(\adder_4bit_13.s<1> ),    .cin(\adder_5bit_6.c<0> ),    .cout(\adder_5bit_6.c<1> ),    .s(\adder_5bit_6.s<1> )
  );
  full_adder \adder_5bit_6.fa_2  (    .a(\adder_4bit_12.s<2> ),    .b(\adder_4bit_13.s<2> ),    .cin(\adder_5bit_6.c<1> ),    .cout(\adder_5bit_6.c<2> ),    .s(\adder_5bit_6.s<2> )
  );
  full_adder \adder_5bit_6.fa_3  (    .a(\adder_4bit_12.s<3> ),    .b(\adder_4bit_13.s<3> ),    .cin(\adder_5bit_6.c<2> ),    .cout(\adder_5bit_6.c<3> ),    .s(\adder_5bit_6.s<3> )
  );
  full_adder \adder_5bit_6.fa_4  (    .a(\adder_4bit_12.s<4> ),    .b(\adder_4bit_13.s<4> ),    .cin(\adder_5bit_6.c<3> ),    .cout(\adder_5bit_6.c<4> ),    .s(\adder_5bit_6.s<4> )
  );
  adder_sign_extension \adder_5bit_6.fa_5  (    .a(\adder_4bit_12.s<4> ),    .b(\adder_4bit_13.s<4> ),    .cin(\adder_5bit_6.c<4> ),    .s(\adder_5bit_6.s<5> ),    .sign(sign_weight)
  );
  half_adder \adder_5bit_6.ha_0  (    .a(\adder_4bit_12.s<0> ),    .b(\adder_4bit_13.s<0> ),    .cout(\adder_5bit_6.c<0> ),    .s(\adder_5bit_6.s<0> )
  );
  full_adder \adder_5bit_7.fa_1  (    .a(\adder_4bit_14.s<1> ),    .b(\adder_4bit_15.s<1> ),    .cin(\adder_5bit_7.c<0> ),    .cout(\adder_5bit_7.c<1> ),    .s(\adder_5bit_7.s<1> )
  );
  full_adder \adder_5bit_7.fa_2  (    .a(\adder_4bit_14.s<2> ),    .b(\adder_4bit_15.s<2> ),    .cin(\adder_5bit_7.c<1> ),    .cout(\adder_5bit_7.c<2> ),    .s(\adder_5bit_7.s<2> )
  );
  full_adder \adder_5bit_7.fa_3  (    .a(\adder_4bit_14.s<3> ),    .b(\adder_4bit_15.s<3> ),    .cin(\adder_5bit_7.c<2> ),    .cout(\adder_5bit_7.c<3> ),    .s(\adder_5bit_7.s<3> )
  );
  full_adder \adder_5bit_7.fa_4  (    .a(\adder_4bit_14.s<4> ),    .b(\adder_4bit_15.s<4> ),    .cin(\adder_5bit_7.c<3> ),    .cout(\adder_5bit_7.c<4> ),    .s(\adder_5bit_7.s<4> )
  );
  adder_sign_extension \adder_5bit_7.fa_5  (    .a(\adder_4bit_14.s<4> ),    .b(\adder_4bit_15.s<4> ),    .cin(\adder_5bit_7.c<4> ),    .s(\adder_5bit_7.s<5> ),    .sign(sign_weight)
  );
  half_adder \adder_5bit_7.ha_0  (    .a(\adder_4bit_14.s<0> ),    .b(\adder_4bit_15.s<0> ),    .cout(\adder_5bit_7.c<0> ),    .s(\adder_5bit_7.s<0> )
  );
  full_adder \adder_5bit_8.fa_1  (    .a(\adder_4bit_16.s<1> ),    .b(\adder_4bit_17.s<1> ),    .cin(\adder_5bit_8.c<0> ),    .cout(\adder_5bit_8.c<1> ),    .s(\adder_5bit_8.s<1> )
  );
  full_adder \adder_5bit_8.fa_2  (    .a(\adder_4bit_16.s<2> ),    .b(\adder_4bit_17.s<2> ),    .cin(\adder_5bit_8.c<1> ),    .cout(\adder_5bit_8.c<2> ),    .s(\adder_5bit_8.s<2> )
  );
  full_adder \adder_5bit_8.fa_3  (    .a(\adder_4bit_16.s<3> ),    .b(\adder_4bit_17.s<3> ),    .cin(\adder_5bit_8.c<2> ),    .cout(\adder_5bit_8.c<3> ),    .s(\adder_5bit_8.s<3> )
  );
  full_adder \adder_5bit_8.fa_4  (    .a(\adder_4bit_16.s<4> ),    .b(\adder_4bit_17.s<4> ),    .cin(\adder_5bit_8.c<3> ),    .cout(\adder_5bit_8.c<4> ),    .s(\adder_5bit_8.s<4> )
  );
  adder_sign_extension \adder_5bit_8.fa_5  (    .a(\adder_4bit_16.s<4> ),    .b(\adder_4bit_17.s<4> ),    .cin(\adder_5bit_8.c<4> ),    .s(\adder_5bit_8.s<5> ),    .sign(sign_weight)
  );
  half_adder \adder_5bit_8.ha_0  (    .a(\adder_4bit_16.s<0> ),    .b(\adder_4bit_17.s<0> ),    .cout(\adder_5bit_8.c<0> ),    .s(\adder_5bit_8.s<0> )
  );
  full_adder \adder_5bit_9.fa_1  (    .a(\adder_4bit_18.s<1> ),    .b(\adder_4bit_19.s<1> ),    .cin(\adder_5bit_9.c<0> ),    .cout(\adder_5bit_9.c<1> ),    .s(\adder_5bit_9.s<1> )
  );
  full_adder \adder_5bit_9.fa_2  (    .a(\adder_4bit_18.s<2> ),    .b(\adder_4bit_19.s<2> ),    .cin(\adder_5bit_9.c<1> ),    .cout(\adder_5bit_9.c<2> ),    .s(\adder_5bit_9.s<2> )
  );
  full_adder \adder_5bit_9.fa_3  (    .a(\adder_4bit_18.s<3> ),    .b(\adder_4bit_19.s<3> ),    .cin(\adder_5bit_9.c<2> ),    .cout(\adder_5bit_9.c<3> ),    .s(\adder_5bit_9.s<3> )
  );
  full_adder \adder_5bit_9.fa_4  (    .a(\adder_4bit_18.s<4> ),    .b(\adder_4bit_19.s<4> ),    .cin(\adder_5bit_9.c<3> ),    .cout(\adder_5bit_9.c<4> ),    .s(\adder_5bit_9.s<4> )
  );
  adder_sign_extension \adder_5bit_9.fa_5  (    .a(\adder_4bit_18.s<4> ),    .b(\adder_4bit_19.s<4> ),    .cin(\adder_5bit_9.c<4> ),    .s(\adder_5bit_9.s<5> ),    .sign(sign_weight)
  );
  half_adder \adder_5bit_9.ha_0  (    .a(\adder_4bit_18.s<0> ),    .b(\adder_4bit_19.s<0> ),    .cout(\adder_5bit_9.c<0> ),    .s(\adder_5bit_9.s<0> )
  );
  full_adder \adder_6bit_0.fa_1  (    .a(\adder_5bit_0.s<1> ),    .b(\adder_5bit_1.s<1> ),    .cin(\adder_6bit_0.c<0> ),    .cout(\adder_6bit_0.c<1> ),    .s(\adder_6bit_0.s<1> )
  );
  full_adder \adder_6bit_0.fa_2  (    .a(\adder_5bit_0.s<2> ),    .b(\adder_5bit_1.s<2> ),    .cin(\adder_6bit_0.c<1> ),    .cout(\adder_6bit_0.c<2> ),    .s(\adder_6bit_0.s<2> )
  );
  full_adder \adder_6bit_0.fa_3  (    .a(\adder_5bit_0.s<3> ),    .b(\adder_5bit_1.s<3> ),    .cin(\adder_6bit_0.c<2> ),    .cout(\adder_6bit_0.c<3> ),    .s(\adder_6bit_0.s<3> )
  );
  full_adder \adder_6bit_0.fa_4  (    .a(\adder_5bit_0.s<4> ),    .b(\adder_5bit_1.s<4> ),    .cin(\adder_6bit_0.c<3> ),    .cout(\adder_6bit_0.c<4> ),    .s(\adder_6bit_0.s<4> )
  );
  full_adder \adder_6bit_0.fa_5  (    .a(\adder_5bit_0.s<5> ),    .b(\adder_5bit_1.s<5> ),    .cin(\adder_6bit_0.c<4> ),    .cout(\adder_6bit_0.c<5> ),    .s(\adder_6bit_0.s<5> )
  );
  adder_sign_extension \adder_6bit_0.fa_6  (    .a(\adder_5bit_0.s<5> ),    .b(\adder_5bit_1.s<5> ),    .cin(\adder_6bit_0.c<5> ),    .s(\adder_6bit_0.s<6> ),    .sign(sign_weight)
  );
  half_adder \adder_6bit_0.ha_0  (    .a(\adder_5bit_0.s<0> ),    .b(\adder_5bit_1.s<0> ),    .cout(\adder_6bit_0.c<0> ),    .s(\adder_6bit_0.s<0> )
  );
  full_adder \adder_6bit_1.fa_1  (    .a(\adder_5bit_2.s<1> ),    .b(\adder_5bit_3.s<1> ),    .cin(\adder_6bit_1.c<0> ),    .cout(\adder_6bit_1.c<1> ),    .s(\adder_6bit_1.s<1> )
  );
  full_adder \adder_6bit_1.fa_2  (    .a(\adder_5bit_2.s<2> ),    .b(\adder_5bit_3.s<2> ),    .cin(\adder_6bit_1.c<1> ),    .cout(\adder_6bit_1.c<2> ),    .s(\adder_6bit_1.s<2> )
  );
  full_adder \adder_6bit_1.fa_3  (    .a(\adder_5bit_2.s<3> ),    .b(\adder_5bit_3.s<3> ),    .cin(\adder_6bit_1.c<2> ),    .cout(\adder_6bit_1.c<3> ),    .s(\adder_6bit_1.s<3> )
  );
  full_adder \adder_6bit_1.fa_4  (    .a(\adder_5bit_2.s<4> ),    .b(\adder_5bit_3.s<4> ),    .cin(\adder_6bit_1.c<3> ),    .cout(\adder_6bit_1.c<4> ),    .s(\adder_6bit_1.s<4> )
  );
  full_adder \adder_6bit_1.fa_5  (    .a(\adder_5bit_2.s<5> ),    .b(\adder_5bit_3.s<5> ),    .cin(\adder_6bit_1.c<4> ),    .cout(\adder_6bit_1.c<5> ),    .s(\adder_6bit_1.s<5> )
  );
  adder_sign_extension \adder_6bit_1.fa_6  (    .a(\adder_5bit_2.s<5> ),    .b(\adder_5bit_3.s<5> ),    .cin(\adder_6bit_1.c<5> ),    .s(\adder_6bit_1.s<6> ),    .sign(sign_weight)
  );
  half_adder \adder_6bit_1.ha_0  (    .a(\adder_5bit_2.s<0> ),    .b(\adder_5bit_3.s<0> ),    .cout(\adder_6bit_1.c<0> ),    .s(\adder_6bit_1.s<0> )
  );
  full_adder \adder_6bit_2.fa_1  (    .a(\adder_5bit_4.s<1> ),    .b(\adder_5bit_5.s<1> ),    .cin(\adder_6bit_2.c<0> ),    .cout(\adder_6bit_2.c<1> ),    .s(\adder_6bit_2.s<1> )
  );
  full_adder \adder_6bit_2.fa_2  (    .a(\adder_5bit_4.s<2> ),    .b(\adder_5bit_5.s<2> ),    .cin(\adder_6bit_2.c<1> ),    .cout(\adder_6bit_2.c<2> ),    .s(\adder_6bit_2.s<2> )
  );
  full_adder \adder_6bit_2.fa_3  (    .a(\adder_5bit_4.s<3> ),    .b(\adder_5bit_5.s<3> ),    .cin(\adder_6bit_2.c<2> ),    .cout(\adder_6bit_2.c<3> ),    .s(\adder_6bit_2.s<3> )
  );
  full_adder \adder_6bit_2.fa_4  (    .a(\adder_5bit_4.s<4> ),    .b(\adder_5bit_5.s<4> ),    .cin(\adder_6bit_2.c<3> ),    .cout(\adder_6bit_2.c<4> ),    .s(\adder_6bit_2.s<4> )
  );
  full_adder \adder_6bit_2.fa_5  (    .a(\adder_5bit_4.s<5> ),    .b(\adder_5bit_5.s<5> ),    .cin(\adder_6bit_2.c<4> ),    .cout(\adder_6bit_2.c<5> ),    .s(\adder_6bit_2.s<5> )
  );
  adder_sign_extension \adder_6bit_2.fa_6  (    .a(\adder_5bit_4.s<5> ),    .b(\adder_5bit_5.s<5> ),    .cin(\adder_6bit_2.c<5> ),    .s(\adder_6bit_2.s<6> ),    .sign(sign_weight)
  );
  half_adder \adder_6bit_2.ha_0  (    .a(\adder_5bit_4.s<0> ),    .b(\adder_5bit_5.s<0> ),    .cout(\adder_6bit_2.c<0> ),    .s(\adder_6bit_2.s<0> )
  );
  full_adder \adder_6bit_3.fa_1  (    .a(\adder_5bit_6.s<1> ),    .b(\adder_5bit_7.s<1> ),    .cin(\adder_6bit_3.c<0> ),    .cout(\adder_6bit_3.c<1> ),    .s(\adder_6bit_3.s<1> )
  );
  full_adder \adder_6bit_3.fa_2  (    .a(\adder_5bit_6.s<2> ),    .b(\adder_5bit_7.s<2> ),    .cin(\adder_6bit_3.c<1> ),    .cout(\adder_6bit_3.c<2> ),    .s(\adder_6bit_3.s<2> )
  );
  full_adder \adder_6bit_3.fa_3  (    .a(\adder_5bit_6.s<3> ),    .b(\adder_5bit_7.s<3> ),    .cin(\adder_6bit_3.c<2> ),    .cout(\adder_6bit_3.c<3> ),    .s(\adder_6bit_3.s<3> )
  );
  full_adder \adder_6bit_3.fa_4  (    .a(\adder_5bit_6.s<4> ),    .b(\adder_5bit_7.s<4> ),    .cin(\adder_6bit_3.c<3> ),    .cout(\adder_6bit_3.c<4> ),    .s(\adder_6bit_3.s<4> )
  );
  full_adder \adder_6bit_3.fa_5  (    .a(\adder_5bit_6.s<5> ),    .b(\adder_5bit_7.s<5> ),    .cin(\adder_6bit_3.c<4> ),    .cout(\adder_6bit_3.c<5> ),    .s(\adder_6bit_3.s<5> )
  );
  adder_sign_extension \adder_6bit_3.fa_6  (    .a(\adder_5bit_6.s<5> ),    .b(\adder_5bit_7.s<5> ),    .cin(\adder_6bit_3.c<5> ),    .s(\adder_6bit_3.s<6> ),    .sign(sign_weight)
  );
  half_adder \adder_6bit_3.ha_0  (    .a(\adder_5bit_6.s<0> ),    .b(\adder_5bit_7.s<0> ),    .cout(\adder_6bit_3.c<0> ),    .s(\adder_6bit_3.s<0> )
  );
  full_adder \adder_6bit_4.fa_1  (    .a(\adder_5bit_8.s<1> ),    .b(\adder_5bit_9.s<1> ),    .cin(\adder_6bit_4.c<0> ),    .cout(\adder_6bit_4.c<1> ),    .s(\adder_6bit_4.s<1> )
  );
  full_adder \adder_6bit_4.fa_2  (    .a(\adder_5bit_8.s<2> ),    .b(\adder_5bit_9.s<2> ),    .cin(\adder_6bit_4.c<1> ),    .cout(\adder_6bit_4.c<2> ),    .s(\adder_6bit_4.s<2> )
  );
  full_adder \adder_6bit_4.fa_3  (    .a(\adder_5bit_8.s<3> ),    .b(\adder_5bit_9.s<3> ),    .cin(\adder_6bit_4.c<2> ),    .cout(\adder_6bit_4.c<3> ),    .s(\adder_6bit_4.s<3> )
  );
  full_adder \adder_6bit_4.fa_4  (    .a(\adder_5bit_8.s<4> ),    .b(\adder_5bit_9.s<4> ),    .cin(\adder_6bit_4.c<3> ),    .cout(\adder_6bit_4.c<4> ),    .s(\adder_6bit_4.s<4> )
  );
  full_adder \adder_6bit_4.fa_5  (    .a(\adder_5bit_8.s<5> ),    .b(\adder_5bit_9.s<5> ),    .cin(\adder_6bit_4.c<4> ),    .cout(\adder_6bit_4.c<5> ),    .s(\adder_6bit_4.s<5> )
  );
  adder_sign_extension \adder_6bit_4.fa_6  (    .a(\adder_5bit_8.s<5> ),    .b(\adder_5bit_9.s<5> ),    .cin(\adder_6bit_4.c<5> ),    .s(\adder_6bit_4.s<6> ),    .sign(sign_weight)
  );
  half_adder \adder_6bit_4.ha_0  (    .a(\adder_5bit_8.s<0> ),    .b(\adder_5bit_9.s<0> ),    .cout(\adder_6bit_4.c<0> ),    .s(\adder_6bit_4.s<0> )
  );
  full_adder \adder_6bit_5.fa_1  (    .a(\adder_5bit_10.s<1> ),    .b(\adder_5bit_11.s<1> ),    .cin(\adder_6bit_5.c<0> ),    .cout(\adder_6bit_5.c<1> ),    .s(\adder_6bit_5.s<1> )
  );
  full_adder \adder_6bit_5.fa_2  (    .a(\adder_5bit_10.s<2> ),    .b(\adder_5bit_11.s<2> ),    .cin(\adder_6bit_5.c<1> ),    .cout(\adder_6bit_5.c<2> ),    .s(\adder_6bit_5.s<2> )
  );
  full_adder \adder_6bit_5.fa_3  (    .a(\adder_5bit_10.s<3> ),    .b(\adder_5bit_11.s<3> ),    .cin(\adder_6bit_5.c<2> ),    .cout(\adder_6bit_5.c<3> ),    .s(\adder_6bit_5.s<3> )
  );
  full_adder \adder_6bit_5.fa_4  (    .a(\adder_5bit_10.s<4> ),    .b(\adder_5bit_11.s<4> ),    .cin(\adder_6bit_5.c<3> ),    .cout(\adder_6bit_5.c<4> ),    .s(\adder_6bit_5.s<4> )
  );
  full_adder \adder_6bit_5.fa_5  (    .a(\adder_5bit_10.s<5> ),    .b(\adder_5bit_11.s<5> ),    .cin(\adder_6bit_5.c<4> ),    .cout(\adder_6bit_5.c<5> ),    .s(\adder_6bit_5.s<5> )
  );
  adder_sign_extension \adder_6bit_5.fa_6  (    .a(\adder_5bit_10.s<5> ),    .b(\adder_5bit_11.s<5> ),    .cin(\adder_6bit_5.c<5> ),    .s(\adder_6bit_5.s<6> ),    .sign(sign_weight)
  );
  half_adder \adder_6bit_5.ha_0  (    .a(\adder_5bit_10.s<0> ),    .b(\adder_5bit_11.s<0> ),    .cout(\adder_6bit_5.c<0> ),    .s(\adder_6bit_5.s<0> )
  );
  full_adder \adder_6bit_6.fa_1  (    .a(\adder_5bit_12.s<1> ),    .b(\adder_5bit_13.s<1> ),    .cin(\adder_6bit_6.c<0> ),    .cout(\adder_6bit_6.c<1> ),    .s(\adder_6bit_6.s<1> )
  );
  full_adder \adder_6bit_6.fa_2  (    .a(\adder_5bit_12.s<2> ),    .b(\adder_5bit_13.s<2> ),    .cin(\adder_6bit_6.c<1> ),    .cout(\adder_6bit_6.c<2> ),    .s(\adder_6bit_6.s<2> )
  );
  full_adder \adder_6bit_6.fa_3  (    .a(\adder_5bit_12.s<3> ),    .b(\adder_5bit_13.s<3> ),    .cin(\adder_6bit_6.c<2> ),    .cout(\adder_6bit_6.c<3> ),    .s(\adder_6bit_6.s<3> )
  );
  full_adder \adder_6bit_6.fa_4  (    .a(\adder_5bit_12.s<4> ),    .b(\adder_5bit_13.s<4> ),    .cin(\adder_6bit_6.c<3> ),    .cout(\adder_6bit_6.c<4> ),    .s(\adder_6bit_6.s<4> )
  );
  full_adder \adder_6bit_6.fa_5  (    .a(\adder_5bit_12.s<5> ),    .b(\adder_5bit_13.s<5> ),    .cin(\adder_6bit_6.c<4> ),    .cout(\adder_6bit_6.c<5> ),    .s(\adder_6bit_6.s<5> )
  );
  adder_sign_extension \adder_6bit_6.fa_6  (    .a(\adder_5bit_12.s<5> ),    .b(\adder_5bit_13.s<5> ),    .cin(\adder_6bit_6.c<5> ),    .s(\adder_6bit_6.s<6> ),    .sign(sign_weight)
  );
  half_adder \adder_6bit_6.ha_0  (    .a(\adder_5bit_12.s<0> ),    .b(\adder_5bit_13.s<0> ),    .cout(\adder_6bit_6.c<0> ),    .s(\adder_6bit_6.s<0> )
  );
  full_adder \adder_6bit_7.fa_1  (    .a(\adder_5bit_14.s<1> ),    .b(\adder_5bit_15.s<1> ),    .cin(\adder_6bit_7.c<0> ),    .cout(\adder_6bit_7.c<1> ),    .s(\adder_6bit_7.s<1> )
  );
  full_adder \adder_6bit_7.fa_2  (    .a(\adder_5bit_14.s<2> ),    .b(\adder_5bit_15.s<2> ),    .cin(\adder_6bit_7.c<1> ),    .cout(\adder_6bit_7.c<2> ),    .s(\adder_6bit_7.s<2> )
  );
  full_adder \adder_6bit_7.fa_3  (    .a(\adder_5bit_14.s<3> ),    .b(\adder_5bit_15.s<3> ),    .cin(\adder_6bit_7.c<2> ),    .cout(\adder_6bit_7.c<3> ),    .s(\adder_6bit_7.s<3> )
  );
  full_adder \adder_6bit_7.fa_4  (    .a(\adder_5bit_14.s<4> ),    .b(\adder_5bit_15.s<4> ),    .cin(\adder_6bit_7.c<3> ),    .cout(\adder_6bit_7.c<4> ),    .s(\adder_6bit_7.s<4> )
  );
  full_adder \adder_6bit_7.fa_5  (    .a(\adder_5bit_14.s<5> ),    .b(\adder_5bit_15.s<5> ),    .cin(\adder_6bit_7.c<4> ),    .cout(\adder_6bit_7.c<5> ),    .s(\adder_6bit_7.s<5> )
  );
  adder_sign_extension \adder_6bit_7.fa_6  (    .a(\adder_5bit_14.s<5> ),    .b(\adder_5bit_15.s<5> ),    .cin(\adder_6bit_7.c<5> ),    .s(\adder_6bit_7.s<6> ),    .sign(sign_weight)
  );
  half_adder \adder_6bit_7.ha_0  (    .a(\adder_5bit_14.s<0> ),    .b(\adder_5bit_15.s<0> ),    .cout(\adder_6bit_7.c<0> ),    .s(\adder_6bit_7.s<0> )
  );
  full_adder \adder_7bit_0.fa_1  (    .a(\adder_6bit_0.s<1> ),    .b(\adder_6bit_1.s<1> ),    .cin(\adder_7bit_0.c<0> ),    .cout(\adder_7bit_0.c<1> ),    .s(\adder_7bit_0.s<1> )
  );
  full_adder \adder_7bit_0.fa_2  (    .a(\adder_6bit_0.s<2> ),    .b(\adder_6bit_1.s<2> ),    .cin(\adder_7bit_0.c<1> ),    .cout(\adder_7bit_0.c<2> ),    .s(\adder_7bit_0.s<2> )
  );
  full_adder \adder_7bit_0.fa_3  (    .a(\adder_6bit_0.s<3> ),    .b(\adder_6bit_1.s<3> ),    .cin(\adder_7bit_0.c<2> ),    .cout(\adder_7bit_0.c<3> ),    .s(\adder_7bit_0.s<3> )
  );
  full_adder \adder_7bit_0.fa_4  (    .a(\adder_6bit_0.s<4> ),    .b(\adder_6bit_1.s<4> ),    .cin(\adder_7bit_0.c<3> ),    .cout(\adder_7bit_0.c<4> ),    .s(\adder_7bit_0.s<4> )
  );
  full_adder \adder_7bit_0.fa_5  (    .a(\adder_6bit_0.s<5> ),    .b(\adder_6bit_1.s<5> ),    .cin(\adder_7bit_0.c<4> ),    .cout(\adder_7bit_0.c<5> ),    .s(\adder_7bit_0.s<5> )
  );
  full_adder \adder_7bit_0.fa_6  (    .a(\adder_6bit_0.s<6> ),    .b(\adder_6bit_1.s<6> ),    .cin(\adder_7bit_0.c<5> ),    .cout(\adder_7bit_0.c<6> ),    .s(\adder_7bit_0.s<6> )
  );
  adder_sign_extension \adder_7bit_0.fa_7  (    .a(\adder_6bit_0.s<6> ),    .b(\adder_6bit_1.s<6> ),    .cin(\adder_7bit_0.c<6> ),    .s(\adder_7bit_0.s<7> ),    .sign(sign_weight)
  );
  half_adder \adder_7bit_0.ha_0  (    .a(\adder_6bit_0.s<0> ),    .b(\adder_6bit_1.s<0> ),    .cout(\adder_7bit_0.c<0> ),    .s(\adder_7bit_0.s<0> )
  );
  full_adder \adder_7bit_1.fa_1  (    .a(\adder_6bit_2.s<1> ),    .b(\adder_6bit_3.s<1> ),    .cin(\adder_7bit_1.c<0> ),    .cout(\adder_7bit_1.c<1> ),    .s(\adder_7bit_1.s<1> )
  );
  full_adder \adder_7bit_1.fa_2  (    .a(\adder_6bit_2.s<2> ),    .b(\adder_6bit_3.s<2> ),    .cin(\adder_7bit_1.c<1> ),    .cout(\adder_7bit_1.c<2> ),    .s(\adder_7bit_1.s<2> )
  );
  full_adder \adder_7bit_1.fa_3  (    .a(\adder_6bit_2.s<3> ),    .b(\adder_6bit_3.s<3> ),    .cin(\adder_7bit_1.c<2> ),    .cout(\adder_7bit_1.c<3> ),    .s(\adder_7bit_1.s<3> )
  );
  full_adder \adder_7bit_1.fa_4  (    .a(\adder_6bit_2.s<4> ),    .b(\adder_6bit_3.s<4> ),    .cin(\adder_7bit_1.c<3> ),    .cout(\adder_7bit_1.c<4> ),    .s(\adder_7bit_1.s<4> )
  );
  full_adder \adder_7bit_1.fa_5  (    .a(\adder_6bit_2.s<5> ),    .b(\adder_6bit_3.s<5> ),    .cin(\adder_7bit_1.c<4> ),    .cout(\adder_7bit_1.c<5> ),    .s(\adder_7bit_1.s<5> )
  );
  full_adder \adder_7bit_1.fa_6  (    .a(\adder_6bit_2.s<6> ),    .b(\adder_6bit_3.s<6> ),    .cin(\adder_7bit_1.c<5> ),    .cout(\adder_7bit_1.c<6> ),    .s(\adder_7bit_1.s<6> )
  );
  adder_sign_extension \adder_7bit_1.fa_7  (    .a(\adder_6bit_2.s<6> ),    .b(\adder_6bit_3.s<6> ),    .cin(\adder_7bit_1.c<6> ),    .s(\adder_7bit_1.s<7> ),    .sign(sign_weight)
  );
  half_adder \adder_7bit_1.ha_0  (    .a(\adder_6bit_2.s<0> ),    .b(\adder_6bit_3.s<0> ),    .cout(\adder_7bit_1.c<0> ),    .s(\adder_7bit_1.s<0> )
  );
  full_adder \adder_7bit_2.fa_1  (    .a(\adder_6bit_4.s<1> ),    .b(\adder_6bit_5.s<1> ),    .cin(\adder_7bit_2.c<0> ),    .cout(\adder_7bit_2.c<1> ),    .s(\adder_7bit_2.s<1> )
  );
  full_adder \adder_7bit_2.fa_2  (    .a(\adder_6bit_4.s<2> ),    .b(\adder_6bit_5.s<2> ),    .cin(\adder_7bit_2.c<1> ),    .cout(\adder_7bit_2.c<2> ),    .s(\adder_7bit_2.s<2> )
  );
  full_adder \adder_7bit_2.fa_3  (    .a(\adder_6bit_4.s<3> ),    .b(\adder_6bit_5.s<3> ),    .cin(\adder_7bit_2.c<2> ),    .cout(\adder_7bit_2.c<3> ),    .s(\adder_7bit_2.s<3> )
  );
  full_adder \adder_7bit_2.fa_4  (    .a(\adder_6bit_4.s<4> ),    .b(\adder_6bit_5.s<4> ),    .cin(\adder_7bit_2.c<3> ),    .cout(\adder_7bit_2.c<4> ),    .s(\adder_7bit_2.s<4> )
  );
  full_adder \adder_7bit_2.fa_5  (    .a(\adder_6bit_4.s<5> ),    .b(\adder_6bit_5.s<5> ),    .cin(\adder_7bit_2.c<4> ),    .cout(\adder_7bit_2.c<5> ),    .s(\adder_7bit_2.s<5> )
  );
  full_adder \adder_7bit_2.fa_6  (    .a(\adder_6bit_4.s<6> ),    .b(\adder_6bit_5.s<6> ),    .cin(\adder_7bit_2.c<5> ),    .cout(\adder_7bit_2.c<6> ),    .s(\adder_7bit_2.s<6> )
  );
  adder_sign_extension \adder_7bit_2.fa_7  (    .a(\adder_6bit_4.s<6> ),    .b(\adder_6bit_5.s<6> ),    .cin(\adder_7bit_2.c<6> ),    .s(\adder_7bit_2.s<7> ),    .sign(sign_weight)
  );
  half_adder \adder_7bit_2.ha_0  (    .a(\adder_6bit_4.s<0> ),    .b(\adder_6bit_5.s<0> ),    .cout(\adder_7bit_2.c<0> ),    .s(\adder_7bit_2.s<0> )
  );
  full_adder \adder_7bit_3.fa_1  (    .a(\adder_6bit_6.s<1> ),    .b(\adder_6bit_7.s<1> ),    .cin(\adder_7bit_3.c<0> ),    .cout(\adder_7bit_3.c<1> ),    .s(\adder_7bit_3.s<1> )
  );
  full_adder \adder_7bit_3.fa_2  (    .a(\adder_6bit_6.s<2> ),    .b(\adder_6bit_7.s<2> ),    .cin(\adder_7bit_3.c<1> ),    .cout(\adder_7bit_3.c<2> ),    .s(\adder_7bit_3.s<2> )
  );
  full_adder \adder_7bit_3.fa_3  (    .a(\adder_6bit_6.s<3> ),    .b(\adder_6bit_7.s<3> ),    .cin(\adder_7bit_3.c<2> ),    .cout(\adder_7bit_3.c<3> ),    .s(\adder_7bit_3.s<3> )
  );
  full_adder \adder_7bit_3.fa_4  (    .a(\adder_6bit_6.s<4> ),    .b(\adder_6bit_7.s<4> ),    .cin(\adder_7bit_3.c<3> ),    .cout(\adder_7bit_3.c<4> ),    .s(\adder_7bit_3.s<4> )
  );
  full_adder \adder_7bit_3.fa_5  (    .a(\adder_6bit_6.s<5> ),    .b(\adder_6bit_7.s<5> ),    .cin(\adder_7bit_3.c<4> ),    .cout(\adder_7bit_3.c<5> ),    .s(\adder_7bit_3.s<5> )
  );
  full_adder \adder_7bit_3.fa_6  (    .a(\adder_6bit_6.s<6> ),    .b(\adder_6bit_7.s<6> ),    .cin(\adder_7bit_3.c<5> ),    .cout(\adder_7bit_3.c<6> ),    .s(\adder_7bit_3.s<6> )
  );
  adder_sign_extension \adder_7bit_3.fa_7  (    .a(\adder_6bit_6.s<6> ),    .b(\adder_6bit_7.s<6> ),    .cin(\adder_7bit_3.c<6> ),    .s(\adder_7bit_3.s<7> ),    .sign(sign_weight)
  );
  half_adder \adder_7bit_3.ha_0  (    .a(\adder_6bit_6.s<0> ),    .b(\adder_6bit_7.s<0> ),    .cout(\adder_7bit_3.c<0> ),    .s(\adder_7bit_3.s<0> )
  );
  full_adder \adder_8bit_0.fa_1  (    .a(\adder_7bit_0.s<1> ),    .b(\adder_7bit_1.s<1> ),    .cin(\adder_8bit_0.c<0> ),    .cout(\adder_8bit_0.c<1> ),    .s(\adder_8bit_0.s<1> )
  );
  full_adder \adder_8bit_0.fa_2  (    .a(\adder_7bit_0.s<2> ),    .b(\adder_7bit_1.s<2> ),    .cin(\adder_8bit_0.c<1> ),    .cout(\adder_8bit_0.c<2> ),    .s(\adder_8bit_0.s<2> )
  );
  full_adder \adder_8bit_0.fa_3  (    .a(\adder_7bit_0.s<3> ),    .b(\adder_7bit_1.s<3> ),    .cin(\adder_8bit_0.c<2> ),    .cout(\adder_8bit_0.c<3> ),    .s(\adder_8bit_0.s<3> )
  );
  full_adder \adder_8bit_0.fa_4  (    .a(\adder_7bit_0.s<4> ),    .b(\adder_7bit_1.s<4> ),    .cin(\adder_8bit_0.c<3> ),    .cout(\adder_8bit_0.c<4> ),    .s(\adder_8bit_0.s<4> )
  );
  full_adder \adder_8bit_0.fa_5  (    .a(\adder_7bit_0.s<5> ),    .b(\adder_7bit_1.s<5> ),    .cin(\adder_8bit_0.c<4> ),    .cout(\adder_8bit_0.c<5> ),    .s(\adder_8bit_0.s<5> )
  );
  full_adder \adder_8bit_0.fa_6  (    .a(\adder_7bit_0.s<6> ),    .b(\adder_7bit_1.s<6> ),    .cin(\adder_8bit_0.c<5> ),    .cout(\adder_8bit_0.c<6> ),    .s(\adder_8bit_0.s<6> )
  );
  full_adder \adder_8bit_0.fa_7  (    .a(\adder_7bit_0.s<7> ),    .b(\adder_7bit_1.s<7> ),    .cin(\adder_8bit_0.c<6> ),    .cout(\adder_8bit_0.c<7> ),    .s(\adder_8bit_0.s<7> )
  );
  adder_sign_extension \adder_8bit_0.fa_8  (    .a(\adder_7bit_0.s<7> ),    .b(\adder_7bit_1.s<7> ),    .cin(\adder_8bit_0.c<7> ),    .s(\adder_8bit_0.s<8> ),    .sign(sign_weight)
  );
  half_adder \adder_8bit_0.ha_0  (    .a(\adder_7bit_0.s<0> ),    .b(\adder_7bit_1.s<0> ),    .cout(\adder_8bit_0.c<0> ),    .s(\adder_8bit_0.s<0> )
  );
  full_adder \adder_8bit_1.fa_1  (    .a(\adder_7bit_2.s<1> ),    .b(\adder_7bit_3.s<1> ),    .cin(\adder_8bit_1.c<0> ),    .cout(\adder_8bit_1.c<1> ),    .s(\adder_8bit_1.s<1> )
  );
  full_adder \adder_8bit_1.fa_2  (    .a(\adder_7bit_2.s<2> ),    .b(\adder_7bit_3.s<2> ),    .cin(\adder_8bit_1.c<1> ),    .cout(\adder_8bit_1.c<2> ),    .s(\adder_8bit_1.s<2> )
  );
  full_adder \adder_8bit_1.fa_3  (    .a(\adder_7bit_2.s<3> ),    .b(\adder_7bit_3.s<3> ),    .cin(\adder_8bit_1.c<2> ),    .cout(\adder_8bit_1.c<3> ),    .s(\adder_8bit_1.s<3> )
  );
  full_adder \adder_8bit_1.fa_4  (    .a(\adder_7bit_2.s<4> ),    .b(\adder_7bit_3.s<4> ),    .cin(\adder_8bit_1.c<3> ),    .cout(\adder_8bit_1.c<4> ),    .s(\adder_8bit_1.s<4> )
  );
  full_adder \adder_8bit_1.fa_5  (    .a(\adder_7bit_2.s<5> ),    .b(\adder_7bit_3.s<5> ),    .cin(\adder_8bit_1.c<4> ),    .cout(\adder_8bit_1.c<5> ),    .s(\adder_8bit_1.s<5> )
  );
  full_adder \adder_8bit_1.fa_6  (    .a(\adder_7bit_2.s<6> ),    .b(\adder_7bit_3.s<6> ),    .cin(\adder_8bit_1.c<5> ),    .cout(\adder_8bit_1.c<6> ),    .s(\adder_8bit_1.s<6> )
  );
  full_adder \adder_8bit_1.fa_7  (    .a(\adder_7bit_2.s<7> ),    .b(\adder_7bit_3.s<7> ),    .cin(\adder_8bit_1.c<6> ),    .cout(\adder_8bit_1.c<7> ),    .s(\adder_8bit_1.s<7> )
  );
  adder_sign_extension \adder_8bit_1.fa_8  (    .a(\adder_7bit_2.s<7> ),    .b(\adder_7bit_3.s<7> ),    .cin(\adder_8bit_1.c<7> ),    .s(\adder_8bit_1.s<8> ),    .sign(sign_weight)
  );
  half_adder \adder_8bit_1.ha_0  (    .a(\adder_7bit_2.s<0> ),    .b(\adder_7bit_3.s<0> ),    .cout(\adder_8bit_1.c<0> ),    .s(\adder_8bit_1.s<0> )
  );
  full_adder \adder_9bit.fa_1  (    .a(\adder_8bit_0.s<1> ),    .b(\adder_8bit_1.s<1> ),    .cin(\adder_9bit.c<0> ),    .cout(\adder_9bit.c<1> ),    .s(\adder_9bit.s<1> )
  );
  full_adder \adder_9bit.fa_2  (    .a(\adder_8bit_0.s<2> ),    .b(\adder_8bit_1.s<2> ),    .cin(\adder_9bit.c<1> ),    .cout(\adder_9bit.c<2> ),    .s(\adder_9bit.s<2> )
  );
  full_adder \adder_9bit.fa_3  (    .a(\adder_8bit_0.s<3> ),    .b(\adder_8bit_1.s<3> ),    .cin(\adder_9bit.c<2> ),    .cout(\adder_9bit.c<3> ),    .s(\adder_9bit.s<3> )
  );
  full_adder \adder_9bit.fa_4  (    .a(\adder_8bit_0.s<4> ),    .b(\adder_8bit_1.s<4> ),    .cin(\adder_9bit.c<3> ),    .cout(\adder_9bit.c<4> ),    .s(\adder_9bit.s<4> )
  );
  full_adder \adder_9bit.fa_5  (    .a(\adder_8bit_0.s<5> ),    .b(\adder_8bit_1.s<5> ),    .cin(\adder_9bit.c<4> ),    .cout(\adder_9bit.c<5> ),    .s(\adder_9bit.s<5> )
  );
  full_adder \adder_9bit.fa_6  (    .a(\adder_8bit_0.s<6> ),    .b(\adder_8bit_1.s<6> ),    .cin(\adder_9bit.c<5> ),    .cout(\adder_9bit.c<6> ),    .s(\adder_9bit.s<6> )
  );
  full_adder \adder_9bit.fa_7  (    .a(\adder_8bit_0.s<7> ),    .b(\adder_8bit_1.s<7> ),    .cin(\adder_9bit.c<6> ),    .cout(\adder_9bit.c<7> ),    .s(\adder_9bit.s<7> )
  );
  full_adder \adder_9bit.fa_8  (    .a(\adder_8bit_0.s<8> ),    .b(\adder_8bit_1.s<8> ),    .cin(\adder_9bit.c<7> ),    .cout(\adder_9bit.c<8> ),    .s(\adder_9bit.s<8> )
  );
  adder_sign_extension \adder_9bit.fa_9  (    .a(\adder_8bit_0.s<8> ),    .b(\adder_8bit_1.s<8> ),    .cin(\adder_9bit.c<8> ),    .s(\adder_9bit.s<9> ),    .sign(sign_weight)
  );
  half_adder \adder_9bit.ha_0  (    .a(\adder_8bit_0.s<0> ),    .b(\adder_8bit_1.s<0> ),    .cout(\adder_9bit.c<0> ),    .s(\adder_9bit.s<0> )
  );
  assign \adder_7bit_1.a<6>  = \adder_6bit_2.s<6> ;
  assign \adder_7bit_1.a<5>  = \adder_6bit_2.s<5> ;
  assign \adder_7bit_1.a<4>  = \adder_6bit_2.s<4> ;
  assign \adder_7bit_1.a<3>  = \adder_6bit_2.s<3> ;
  assign \adder_7bit_1.a<2>  = \adder_6bit_2.s<2> ;
  assign \adder_7bit_1.a<1>  = \adder_6bit_2.s<1> ;
  assign \adder_7bit_1.a<0>  = \adder_6bit_2.s<0> ;
  assign \adder_7bit_1.b<6>  = \adder_6bit_3.s<6> ;
  assign \adder_7bit_1.b<5>  = \adder_6bit_3.s<5> ;
  assign \adder_7bit_1.b<4>  = \adder_6bit_3.s<4> ;
  assign \adder_7bit_1.b<3>  = \adder_6bit_3.s<3> ;
  assign \adder_7bit_1.b<2>  = \adder_6bit_3.s<2> ;
  assign \adder_7bit_1.b<1>  = \adder_6bit_3.s<1> ;
  assign \adder_7bit_1.b<0>  = \adder_6bit_3.s<0> ;
  assign \adder_7bit_0.a<6>  = \adder_6bit_0.s<6> ;
  assign \adder_7bit_0.a<5>  = \adder_6bit_0.s<5> ;
  assign \adder_7bit_0.a<4>  = \adder_6bit_0.s<4> ;
  assign \adder_7bit_0.a<3>  = \adder_6bit_0.s<3> ;
  assign \adder_7bit_0.a<2>  = \adder_6bit_0.s<2> ;
  assign \adder_7bit_0.a<1>  = \adder_6bit_0.s<1> ;
  assign \adder_7bit_0.a<0>  = \adder_6bit_0.s<0> ;
  assign \adder_7bit_0.b<6>  = \adder_6bit_1.s<6> ;
  assign \adder_7bit_0.b<5>  = \adder_6bit_1.s<5> ;
  assign \adder_7bit_0.b<4>  = \adder_6bit_1.s<4> ;
  assign \adder_7bit_0.b<3>  = \adder_6bit_1.s<3> ;
  assign \adder_7bit_0.b<2>  = \adder_6bit_1.s<2> ;
  assign \adder_7bit_0.b<1>  = \adder_6bit_1.s<1> ;
  assign \adder_7bit_0.b<0>  = \adder_6bit_1.s<0> ;
  assign \adder_6bit_7.a<5>  = \adder_5bit_14.s<5> ;
  assign \adder_6bit_7.a<4>  = \adder_5bit_14.s<4> ;
  assign \adder_6bit_7.a<3>  = \adder_5bit_14.s<3> ;
  assign \adder_6bit_7.a<2>  = \adder_5bit_14.s<2> ;
  assign \adder_6bit_7.a<1>  = \adder_5bit_14.s<1> ;
  assign \adder_6bit_7.a<0>  = \adder_5bit_14.s<0> ;
  assign \adder_6bit_6.a<5>  = \adder_5bit_12.s<5> ;
  assign \adder_6bit_6.a<4>  = \adder_5bit_12.s<4> ;
  assign \adder_6bit_6.a<3>  = \adder_5bit_12.s<3> ;
  assign \adder_6bit_6.a<2>  = \adder_5bit_12.s<2> ;
  assign \adder_6bit_6.a<1>  = \adder_5bit_12.s<1> ;
  assign \adder_6bit_6.a<0>  = \adder_5bit_12.s<0> ;
  assign \adder_6bit_6.b<5>  = \adder_5bit_13.s<5> ;
  assign \adder_6bit_6.b<4>  = \adder_5bit_13.s<4> ;
  assign \adder_6bit_6.b<3>  = \adder_5bit_13.s<3> ;
  assign \adder_6bit_6.b<2>  = \adder_5bit_13.s<2> ;
  assign \adder_6bit_6.b<1>  = \adder_5bit_13.s<1> ;
  assign \adder_6bit_6.b<0>  = \adder_5bit_13.s<0> ;
  assign \adder_6bit_4.a<5>  = \adder_5bit_8.s<5> ;
  assign \adder_6bit_4.a<4>  = \adder_5bit_8.s<4> ;
  assign \adder_6bit_4.a<3>  = \adder_5bit_8.s<3> ;
  assign \adder_6bit_4.a<2>  = \adder_5bit_8.s<2> ;
  assign \adder_6bit_4.a<1>  = \adder_5bit_8.s<1> ;
  assign \adder_6bit_4.a<0>  = \adder_5bit_8.s<0> ;
  assign \adder_6bit_4.b<5>  = \adder_5bit_9.s<5> ;
  assign \adder_6bit_4.b<4>  = \adder_5bit_9.s<4> ;
  assign \adder_6bit_4.b<3>  = \adder_5bit_9.s<3> ;
  assign \adder_6bit_4.b<2>  = \adder_5bit_9.s<2> ;
  assign \adder_6bit_4.b<1>  = \adder_5bit_9.s<1> ;
  assign \adder_6bit_4.b<0>  = \adder_5bit_9.s<0> ;
  assign \adder_6bit_3.a<5>  = \adder_5bit_6.s<5> ;
  assign \adder_6bit_3.a<4>  = \adder_5bit_6.s<4> ;
  assign \adder_6bit_3.a<3>  = \adder_5bit_6.s<3> ;
  assign \adder_6bit_3.a<2>  = \adder_5bit_6.s<2> ;
  assign \adder_6bit_3.a<1>  = \adder_5bit_6.s<1> ;
  assign \adder_6bit_3.a<0>  = \adder_5bit_6.s<0> ;
  assign \adder_6bit_3.b<5>  = \adder_5bit_7.s<5> ;
  assign \adder_6bit_3.b<4>  = \adder_5bit_7.s<4> ;
  assign \adder_6bit_3.b<3>  = \adder_5bit_7.s<3> ;
  assign \adder_6bit_3.b<2>  = \adder_5bit_7.s<2> ;
  assign \adder_6bit_3.b<1>  = \adder_5bit_7.s<1> ;
  assign \adder_6bit_3.b<0>  = \adder_5bit_7.s<0> ;
  assign \adder_6bit_0.a<5>  = \adder_5bit_0.s<5> ;
  assign \adder_6bit_0.a<4>  = \adder_5bit_0.s<4> ;
  assign \adder_6bit_0.a<3>  = \adder_5bit_0.s<3> ;
  assign \adder_6bit_0.a<2>  = \adder_5bit_0.s<2> ;
  assign \adder_6bit_0.a<1>  = \adder_5bit_0.s<1> ;
  assign \adder_6bit_0.a<0>  = \adder_5bit_0.s<0> ;
  assign \adder_5bit_13.a<4>  = \adder_4bit_26.s<4> ;
  assign \adder_5bit_13.a<3>  = \adder_4bit_26.s<3> ;
  assign \adder_5bit_13.a<2>  = \adder_4bit_26.s<2> ;
  assign \adder_5bit_13.a<1>  = \adder_4bit_26.s<1> ;
  assign \adder_5bit_13.a<0>  = \adder_4bit_26.s<0> ;
  assign \adder_5bit_11.a<4>  = \adder_4bit_22.s<4> ;
  assign \adder_5bit_11.a<3>  = \adder_4bit_22.s<3> ;
  assign \adder_5bit_11.a<2>  = \adder_4bit_22.s<2> ;
  assign \adder_5bit_11.a<1>  = \adder_4bit_22.s<1> ;
  assign \adder_5bit_11.a<0>  = \adder_4bit_22.s<0> ;
  assign \adder_5bit_10.a<4>  = \adder_4bit_20.s<4> ;
  assign \adder_5bit_10.a<3>  = \adder_4bit_20.s<3> ;
  assign \adder_5bit_10.a<2>  = \adder_4bit_20.s<2> ;
  assign \adder_5bit_10.a<1>  = \adder_4bit_20.s<1> ;
  assign \adder_5bit_10.a<0>  = \adder_4bit_20.s<0> ;
  assign \adder_5bit_9.a<4>  = \adder_4bit_18.s<4> ;
  assign \adder_5bit_9.a<3>  = \adder_4bit_18.s<3> ;
  assign \adder_5bit_9.a<2>  = \adder_4bit_18.s<2> ;
  assign \adder_5bit_9.a<1>  = \adder_4bit_18.s<1> ;
  assign \adder_5bit_9.a<0>  = \adder_4bit_18.s<0> ;
  assign \adder_5bit_8.a<4>  = \adder_4bit_16.s<4> ;
  assign \adder_5bit_8.a<3>  = \adder_4bit_16.s<3> ;
  assign \adder_5bit_8.a<2>  = \adder_4bit_16.s<2> ;
  assign \adder_5bit_8.a<1>  = \adder_4bit_16.s<1> ;
  assign \adder_5bit_8.a<0>  = \adder_4bit_16.s<0> ;
  assign \adder_5bit_7.a<4>  = \adder_4bit_14.s<4> ;
  assign \adder_5bit_7.a<3>  = \adder_4bit_14.s<3> ;
  assign \adder_5bit_7.a<2>  = \adder_4bit_14.s<2> ;
  assign \adder_5bit_7.a<1>  = \adder_4bit_14.s<1> ;
  assign \adder_5bit_7.a<0>  = \adder_4bit_14.s<0> ;
  assign \adder_5bit_3.a<4>  = \adder_4bit_6.s<4> ;
  assign \adder_5bit_3.a<3>  = \adder_4bit_6.s<3> ;
  assign \adder_5bit_3.a<2>  = \adder_4bit_6.s<2> ;
  assign \adder_5bit_3.a<1>  = \adder_4bit_6.s<1> ;
  assign \adder_5bit_3.a<0>  = \adder_4bit_6.s<0> ;
  assign \adder_5bit_2.a<4>  = \adder_4bit_4.s<4> ;
  assign \adder_5bit_2.a<3>  = \adder_4bit_4.s<3> ;
  assign \adder_5bit_2.a<2>  = \adder_4bit_4.s<2> ;
  assign \adder_5bit_2.a<1>  = \adder_4bit_4.s<1> ;
  assign \adder_5bit_2.a<0>  = \adder_4bit_4.s<0> ;
  assign \adder_5bit_0.a<4>  = \adder_4bit_0.s<4> ;
  assign \adder_5bit_0.a<3>  = \adder_4bit_0.s<3> ;
  assign \adder_5bit_0.a<2>  = \adder_4bit_0.s<2> ;
  assign \adder_5bit_0.a<1>  = \adder_4bit_0.s<1> ;
  assign \adder_5bit_0.a<0>  = \adder_4bit_0.s<0> ;
  assign \adder_5bit_0.b<4>  = \adder_4bit_1.s<4> ;
  assign \adder_5bit_0.b<3>  = \adder_4bit_1.s<3> ;
  assign \adder_5bit_0.b<2>  = \adder_4bit_1.s<2> ;
  assign \adder_5bit_0.b<1>  = \adder_4bit_1.s<1> ;
  assign \adder_5bit_0.b<0>  = \adder_4bit_1.s<0> ;
  assign \adder_4bit_30.a<3>  = \in_60<3> ;
  assign \adder_4bit_30.a<2>  = \in_60<2> ;
  assign \adder_4bit_30.a<1>  = \in_60<1> ;
  assign \adder_4bit_30.a<0>  = \in_60<0> ;
  assign \adder_4bit_29.a<3>  = \in_58<3> ;
  assign \adder_4bit_29.a<2>  = \in_58<2> ;
  assign \adder_4bit_29.a<1>  = \in_58<1> ;
  assign \adder_4bit_29.a<0>  = \in_58<0> ;
  assign \adder_4bit_27.a<3>  = \in_54<3> ;
  assign \adder_4bit_27.a<2>  = \in_54<2> ;
  assign \adder_4bit_27.a<1>  = \in_54<1> ;
  assign \adder_4bit_27.a<0>  = \in_54<0> ;
  assign \adder_4bit_26.a<3>  = \in_52<3> ;
  assign \adder_4bit_26.a<2>  = \in_52<2> ;
  assign \adder_4bit_26.a<1>  = \in_52<1> ;
  assign \adder_4bit_26.a<0>  = \in_52<0> ;
  assign \adder_5bit_1.a<4>  = \adder_4bit_2.s<4> ;
  assign \adder_5bit_1.a<3>  = \adder_4bit_2.s<3> ;
  assign \adder_5bit_1.a<2>  = \adder_4bit_2.s<2> ;
  assign \adder_5bit_1.a<1>  = \adder_4bit_2.s<1> ;
  assign \adder_5bit_1.a<0>  = \adder_4bit_2.s<0> ;
  assign \adder_4bit_25.a<3>  = \in_50<3> ;
  assign \adder_4bit_25.a<2>  = \in_50<2> ;
  assign \adder_4bit_25.a<1>  = \in_50<1> ;
  assign \adder_4bit_25.a<0>  = \in_50<0> ;
  assign \adder_4bit_23.a<3>  = \in_46<3> ;
  assign \adder_4bit_23.a<2>  = \in_46<2> ;
  assign \adder_4bit_23.a<1>  = \in_46<1> ;
  assign \adder_4bit_23.a<0>  = \in_46<0> ;
  assign \adder_4bit_21.a<3>  = \in_42<3> ;
  assign \adder_4bit_21.a<2>  = \in_42<2> ;
  assign \adder_4bit_21.a<1>  = \in_42<1> ;
  assign \adder_4bit_21.a<0>  = \in_42<0> ;
  assign \adder_4bit_20.a<3>  = \in_40<3> ;
  assign \adder_4bit_20.a<2>  = \in_40<2> ;
  assign \adder_4bit_20.a<1>  = \in_40<1> ;
  assign \adder_4bit_20.a<0>  = \in_40<0> ;
  assign \adder_4bit_19.a<3>  = \in_38<3> ;
  assign \adder_4bit_19.a<2>  = \in_38<2> ;
  assign \adder_4bit_19.a<1>  = \in_38<1> ;
  assign \adder_4bit_19.a<0>  = \in_38<0> ;
  assign \adder_4bit_16.a<3>  = \in_32<3> ;
  assign \adder_4bit_16.a<2>  = \in_32<2> ;
  assign \adder_4bit_16.a<1>  = \in_32<1> ;
  assign \adder_4bit_16.a<0>  = \in_32<0> ;
  assign \adder_4bit_15.a<3>  = \in_30<3> ;
  assign \adder_4bit_15.a<2>  = \in_30<2> ;
  assign \adder_4bit_15.a<1>  = \in_30<1> ;
  assign \adder_4bit_15.a<0>  = \in_30<0> ;
  assign \adder_4bit_13.a<3>  = \in_26<3> ;
  assign \adder_4bit_13.a<2>  = \in_26<2> ;
  assign \adder_4bit_13.a<1>  = \in_26<1> ;
  assign \adder_4bit_13.a<0>  = \in_26<0> ;
  assign \adder_4bit_11.a<3>  = \in_22<3> ;
  assign \adder_4bit_11.a<2>  = \in_22<2> ;
  assign \adder_4bit_11.a<1>  = \in_22<1> ;
  assign \adder_4bit_11.a<0>  = \in_22<0> ;
  assign \adder_4bit_10.a<3>  = \in_20<3> ;
  assign \adder_4bit_10.a<2>  = \in_20<2> ;
  assign \adder_4bit_10.a<1>  = \in_20<1> ;
  assign \adder_4bit_10.a<0>  = \in_20<0> ;
  assign \adder_4bit_9.a<3>  = \in_18<3> ;
  assign \adder_4bit_9.a<2>  = \in_18<2> ;
  assign \adder_4bit_9.a<1>  = \in_18<1> ;
  assign \adder_4bit_9.a<0>  = \in_18<0> ;
  assign \adder_4bit_8.a<3>  = \in_16<3> ;
  assign \adder_4bit_8.a<2>  = \in_16<2> ;
  assign \adder_4bit_8.a<1>  = \in_16<1> ;
  assign \adder_4bit_8.a<0>  = \in_16<0> ;
  assign \sum_8bit_1<8>  = \adder_8bit_1.s<8> ;
  assign \sum_8bit_1<7>  = \adder_8bit_1.s<7> ;
  assign \sum_8bit_1<6>  = \adder_8bit_1.s<6> ;
  assign \sum_8bit_1<5>  = \adder_8bit_1.s<5> ;
  assign \sum_8bit_1<4>  = \adder_8bit_1.s<4> ;
  assign \sum_8bit_1<3>  = \adder_8bit_1.s<3> ;
  assign \sum_8bit_1<2>  = \adder_8bit_1.s<2> ;
  assign \sum_8bit_1<1>  = \adder_8bit_1.s<1> ;
  assign \sum_8bit_1<0>  = \adder_8bit_1.s<0> ;
  assign \sum_8bit_0<8>  = \adder_8bit_0.s<8> ;
  assign \sum_8bit_0<7>  = \adder_8bit_0.s<7> ;
  assign \sum_8bit_0<6>  = \adder_8bit_0.s<6> ;
  assign \sum_8bit_0<5>  = \adder_8bit_0.s<5> ;
  assign \sum_8bit_0<4>  = \adder_8bit_0.s<4> ;
  assign \sum_8bit_0<3>  = \adder_8bit_0.s<3> ;
  assign \sum_8bit_0<2>  = \adder_8bit_0.s<2> ;
  assign \sum_8bit_0<1>  = \adder_8bit_0.s<1> ;
  assign \sum_8bit_0<0>  = \adder_8bit_0.s<0> ;
  assign \sum_7bit_3<7>  = \adder_7bit_3.s<7> ;
  assign \sum_7bit_3<6>  = \adder_7bit_3.s<6> ;
  assign \sum_7bit_3<5>  = \adder_7bit_3.s<5> ;
  assign \sum_7bit_3<4>  = \adder_7bit_3.s<4> ;
  assign \sum_7bit_3<3>  = \adder_7bit_3.s<3> ;
  assign \sum_7bit_3<2>  = \adder_7bit_3.s<2> ;
  assign \sum_7bit_3<1>  = \adder_7bit_3.s<1> ;
  assign \sum_7bit_3<0>  = \adder_7bit_3.s<0> ;
  assign \sum_7bit_2<7>  = \adder_7bit_2.s<7> ;
  assign \sum_7bit_2<6>  = \adder_7bit_2.s<6> ;
  assign \sum_7bit_2<5>  = \adder_7bit_2.s<5> ;
  assign \sum_7bit_2<4>  = \adder_7bit_2.s<4> ;
  assign \sum_7bit_2<3>  = \adder_7bit_2.s<3> ;
  assign \sum_7bit_2<2>  = \adder_7bit_2.s<2> ;
  assign \sum_7bit_2<1>  = \adder_7bit_2.s<1> ;
  assign \sum_7bit_2<0>  = \adder_7bit_2.s<0> ;
  assign \sum_7bit_1<7>  = \adder_7bit_1.s<7> ;
  assign \sum_7bit_1<6>  = \adder_7bit_1.s<6> ;
  assign \sum_7bit_1<5>  = \adder_7bit_1.s<5> ;
  assign \sum_7bit_1<4>  = \adder_7bit_1.s<4> ;
  assign \sum_7bit_1<3>  = \adder_7bit_1.s<3> ;
  assign \sum_7bit_1<2>  = \adder_7bit_1.s<2> ;
  assign \sum_7bit_1<1>  = \adder_7bit_1.s<1> ;
  assign \sum_7bit_1<0>  = \adder_7bit_1.s<0> ;
  assign \sum_7bit_0<7>  = \adder_7bit_0.s<7> ;
  assign \sum_7bit_0<6>  = \adder_7bit_0.s<6> ;
  assign \sum_7bit_0<5>  = \adder_7bit_0.s<5> ;
  assign \sum_7bit_0<4>  = \adder_7bit_0.s<4> ;
  assign \sum_7bit_0<3>  = \adder_7bit_0.s<3> ;
  assign \sum_7bit_0<2>  = \adder_7bit_0.s<2> ;
  assign \sum_7bit_0<1>  = \adder_7bit_0.s<1> ;
  assign \sum_7bit_0<0>  = \adder_7bit_0.s<0> ;
  assign \sum_6bit_7<6>  = \adder_6bit_7.s<6> ;
  assign \sum_6bit_7<5>  = \adder_6bit_7.s<5> ;
  assign \sum_6bit_7<4>  = \adder_6bit_7.s<4> ;
  assign \sum_6bit_7<3>  = \adder_6bit_7.s<3> ;
  assign \sum_6bit_7<2>  = \adder_6bit_7.s<2> ;
  assign \sum_6bit_7<1>  = \adder_6bit_7.s<1> ;
  assign \sum_6bit_7<0>  = \adder_6bit_7.s<0> ;
  assign \sum_6bit_6<6>  = \adder_6bit_6.s<6> ;
  assign \sum_6bit_6<5>  = \adder_6bit_6.s<5> ;
  assign \sum_6bit_6<4>  = \adder_6bit_6.s<4> ;
  assign \sum_6bit_6<3>  = \adder_6bit_6.s<3> ;
  assign \sum_6bit_6<2>  = \adder_6bit_6.s<2> ;
  assign \sum_6bit_6<1>  = \adder_6bit_6.s<1> ;
  assign \sum_6bit_6<0>  = \adder_6bit_6.s<0> ;
  assign \sum_6bit_5<6>  = \adder_6bit_5.s<6> ;
  assign \sum_6bit_5<5>  = \adder_6bit_5.s<5> ;
  assign \sum_6bit_5<4>  = \adder_6bit_5.s<4> ;
  assign \sum_6bit_5<3>  = \adder_6bit_5.s<3> ;
  assign \sum_6bit_5<2>  = \adder_6bit_5.s<2> ;
  assign \sum_6bit_5<1>  = \adder_6bit_5.s<1> ;
  assign \sum_6bit_5<0>  = \adder_6bit_5.s<0> ;
  assign \sum_6bit_4<6>  = \adder_6bit_4.s<6> ;
  assign \sum_6bit_4<5>  = \adder_6bit_4.s<5> ;
  assign \sum_6bit_4<4>  = \adder_6bit_4.s<4> ;
  assign \sum_6bit_4<3>  = \adder_6bit_4.s<3> ;
  assign \sum_6bit_4<2>  = \adder_6bit_4.s<2> ;
  assign \sum_6bit_4<1>  = \adder_6bit_4.s<1> ;
  assign \sum_6bit_4<0>  = \adder_6bit_4.s<0> ;
  assign \sum_6bit_3<6>  = \adder_6bit_3.s<6> ;
  assign \sum_6bit_3<5>  = \adder_6bit_3.s<5> ;
  assign \sum_6bit_3<4>  = \adder_6bit_3.s<4> ;
  assign \sum_6bit_3<3>  = \adder_6bit_3.s<3> ;
  assign \sum_6bit_3<2>  = \adder_6bit_3.s<2> ;
  assign \sum_6bit_3<1>  = \adder_6bit_3.s<1> ;
  assign \sum_6bit_3<0>  = \adder_6bit_3.s<0> ;
  assign \sum_6bit_2<6>  = \adder_6bit_2.s<6> ;
  assign \sum_6bit_2<5>  = \adder_6bit_2.s<5> ;
  assign \sum_6bit_2<4>  = \adder_6bit_2.s<4> ;
  assign \sum_6bit_2<3>  = \adder_6bit_2.s<3> ;
  assign \sum_6bit_2<2>  = \adder_6bit_2.s<2> ;
  assign \sum_6bit_2<1>  = \adder_6bit_2.s<1> ;
  assign \sum_6bit_2<0>  = \adder_6bit_2.s<0> ;
  assign \sum_6bit_1<6>  = \adder_6bit_1.s<6> ;
  assign \sum_6bit_1<5>  = \adder_6bit_1.s<5> ;
  assign \sum_6bit_1<4>  = \adder_6bit_1.s<4> ;
  assign \sum_6bit_1<3>  = \adder_6bit_1.s<3> ;
  assign \sum_6bit_1<2>  = \adder_6bit_1.s<2> ;
  assign \sum_6bit_1<1>  = \adder_6bit_1.s<1> ;
  assign \sum_6bit_1<0>  = \adder_6bit_1.s<0> ;
  assign \sum_6bit_0<6>  = \adder_6bit_0.s<6> ;
  assign \sum_6bit_0<5>  = \adder_6bit_0.s<5> ;
  assign \sum_6bit_0<4>  = \adder_6bit_0.s<4> ;
  assign \sum_6bit_0<3>  = \adder_6bit_0.s<3> ;
  assign \sum_6bit_0<2>  = \adder_6bit_0.s<2> ;
  assign \sum_6bit_0<1>  = \adder_6bit_0.s<1> ;
  assign \sum_6bit_0<0>  = \adder_6bit_0.s<0> ;
  assign \sum_5bit_15<5>  = \adder_5bit_15.s<5> ;
  assign \sum_5bit_15<4>  = \adder_5bit_15.s<4> ;
  assign \sum_5bit_15<3>  = \adder_5bit_15.s<3> ;
  assign \sum_5bit_15<2>  = \adder_5bit_15.s<2> ;
  assign \sum_5bit_15<1>  = \adder_5bit_15.s<1> ;
  assign \sum_5bit_15<0>  = \adder_5bit_15.s<0> ;
  assign \sum_5bit_14<5>  = \adder_5bit_14.s<5> ;
  assign \sum_5bit_14<4>  = \adder_5bit_14.s<4> ;
  assign \sum_5bit_14<3>  = \adder_5bit_14.s<3> ;
  assign \sum_5bit_14<2>  = \adder_5bit_14.s<2> ;
  assign \sum_5bit_14<1>  = \adder_5bit_14.s<1> ;
  assign \sum_5bit_14<0>  = \adder_5bit_14.s<0> ;
  assign \sum_5bit_13<5>  = \adder_5bit_13.s<5> ;
  assign \sum_5bit_13<4>  = \adder_5bit_13.s<4> ;
  assign \sum_5bit_13<3>  = \adder_5bit_13.s<3> ;
  assign \sum_5bit_13<2>  = \adder_5bit_13.s<2> ;
  assign \sum_5bit_13<1>  = \adder_5bit_13.s<1> ;
  assign \sum_5bit_13<0>  = \adder_5bit_13.s<0> ;
  assign \sum_5bit_12<5>  = \adder_5bit_12.s<5> ;
  assign \sum_5bit_12<4>  = \adder_5bit_12.s<4> ;
  assign \sum_5bit_12<3>  = \adder_5bit_12.s<3> ;
  assign \sum_5bit_12<2>  = \adder_5bit_12.s<2> ;
  assign \sum_5bit_12<1>  = \adder_5bit_12.s<1> ;
  assign \sum_5bit_12<0>  = \adder_5bit_12.s<0> ;
  assign \sum_5bit_11<5>  = \adder_5bit_11.s<5> ;
  assign \sum_5bit_11<4>  = \adder_5bit_11.s<4> ;
  assign \sum_5bit_11<3>  = \adder_5bit_11.s<3> ;
  assign \sum_5bit_11<2>  = \adder_5bit_11.s<2> ;
  assign \sum_5bit_11<1>  = \adder_5bit_11.s<1> ;
  assign \sum_5bit_11<0>  = \adder_5bit_11.s<0> ;
  assign \sum_5bit_10<5>  = \adder_5bit_10.s<5> ;
  assign \sum_5bit_10<4>  = \adder_5bit_10.s<4> ;
  assign \sum_5bit_10<3>  = \adder_5bit_10.s<3> ;
  assign \sum_5bit_10<2>  = \adder_5bit_10.s<2> ;
  assign \sum_5bit_10<1>  = \adder_5bit_10.s<1> ;
  assign \sum_5bit_10<0>  = \adder_5bit_10.s<0> ;
  assign \sum_5bit_9<5>  = \adder_5bit_9.s<5> ;
  assign \sum_5bit_9<4>  = \adder_5bit_9.s<4> ;
  assign \sum_5bit_9<3>  = \adder_5bit_9.s<3> ;
  assign \sum_5bit_9<2>  = \adder_5bit_9.s<2> ;
  assign \sum_5bit_9<1>  = \adder_5bit_9.s<1> ;
  assign \sum_5bit_9<0>  = \adder_5bit_9.s<0> ;
  assign \sum_5bit_8<5>  = \adder_5bit_8.s<5> ;
  assign \sum_5bit_8<4>  = \adder_5bit_8.s<4> ;
  assign \sum_5bit_8<3>  = \adder_5bit_8.s<3> ;
  assign \sum_5bit_8<2>  = \adder_5bit_8.s<2> ;
  assign \sum_5bit_8<1>  = \adder_5bit_8.s<1> ;
  assign \sum_5bit_8<0>  = \adder_5bit_8.s<0> ;
  assign \sum_5bit_7<5>  = \adder_5bit_7.s<5> ;
  assign \sum_5bit_7<4>  = \adder_5bit_7.s<4> ;
  assign \sum_5bit_7<3>  = \adder_5bit_7.s<3> ;
  assign \sum_5bit_7<2>  = \adder_5bit_7.s<2> ;
  assign \sum_5bit_7<1>  = \adder_5bit_7.s<1> ;
  assign \sum_5bit_7<0>  = \adder_5bit_7.s<0> ;
  assign \sum_5bit_6<5>  = \adder_5bit_6.s<5> ;
  assign \sum_5bit_6<4>  = \adder_5bit_6.s<4> ;
  assign \sum_5bit_6<3>  = \adder_5bit_6.s<3> ;
  assign \sum_5bit_6<2>  = \adder_5bit_6.s<2> ;
  assign \sum_5bit_6<1>  = \adder_5bit_6.s<1> ;
  assign \sum_5bit_6<0>  = \adder_5bit_6.s<0> ;
  assign \sum_5bit_5<5>  = \adder_5bit_5.s<5> ;
  assign \sum_5bit_5<4>  = \adder_5bit_5.s<4> ;
  assign \sum_5bit_5<3>  = \adder_5bit_5.s<3> ;
  assign \sum_5bit_5<2>  = \adder_5bit_5.s<2> ;
  assign \sum_5bit_5<1>  = \adder_5bit_5.s<1> ;
  assign \sum_5bit_5<0>  = \adder_5bit_5.s<0> ;
  assign \sum_5bit_4<5>  = \adder_5bit_4.s<5> ;
  assign \sum_5bit_4<4>  = \adder_5bit_4.s<4> ;
  assign \sum_5bit_4<3>  = \adder_5bit_4.s<3> ;
  assign \sum_5bit_4<2>  = \adder_5bit_4.s<2> ;
  assign \sum_5bit_4<1>  = \adder_5bit_4.s<1> ;
  assign \sum_5bit_4<0>  = \adder_5bit_4.s<0> ;
  assign \sum_5bit_3<5>  = \adder_5bit_3.s<5> ;
  assign \sum_5bit_3<4>  = \adder_5bit_3.s<4> ;
  assign \sum_5bit_3<3>  = \adder_5bit_3.s<3> ;
  assign \sum_5bit_3<2>  = \adder_5bit_3.s<2> ;
  assign \sum_5bit_3<1>  = \adder_5bit_3.s<1> ;
  assign \sum_5bit_3<0>  = \adder_5bit_3.s<0> ;
  assign \sum_5bit_2<5>  = \adder_5bit_2.s<5> ;
  assign \sum_5bit_2<4>  = \adder_5bit_2.s<4> ;
  assign \sum_5bit_2<3>  = \adder_5bit_2.s<3> ;
  assign \sum_5bit_2<2>  = \adder_5bit_2.s<2> ;
  assign \sum_5bit_2<1>  = \adder_5bit_2.s<1> ;
  assign \sum_5bit_2<0>  = \adder_5bit_2.s<0> ;
  assign \sum_5bit_1<5>  = \adder_5bit_1.s<5> ;
  assign \sum_5bit_1<4>  = \adder_5bit_1.s<4> ;
  assign \sum_5bit_1<3>  = \adder_5bit_1.s<3> ;
  assign \sum_5bit_1<2>  = \adder_5bit_1.s<2> ;
  assign \sum_5bit_1<1>  = \adder_5bit_1.s<1> ;
  assign \sum_5bit_1<0>  = \adder_5bit_1.s<0> ;
  assign \sum_5bit_0<5>  = \adder_5bit_0.s<5> ;
  assign \sum_5bit_0<4>  = \adder_5bit_0.s<4> ;
  assign \sum_5bit_0<3>  = \adder_5bit_0.s<3> ;
  assign \sum_5bit_0<2>  = \adder_5bit_0.s<2> ;
  assign \sum_5bit_0<1>  = \adder_5bit_0.s<1> ;
  assign \sum_5bit_0<0>  = \adder_5bit_0.s<0> ;
  assign \sum_4bit_31<4>  = \adder_4bit_31.s<4> ;
  assign \sum_4bit_31<3>  = \adder_4bit_31.s<3> ;
  assign \sum_4bit_31<2>  = \adder_4bit_31.s<2> ;
  assign \sum_4bit_31<1>  = \adder_4bit_31.s<1> ;
  assign \sum_4bit_31<0>  = \adder_4bit_31.s<0> ;
  assign \sum_4bit_30<4>  = \adder_4bit_30.s<4> ;
  assign \sum_4bit_30<3>  = \adder_4bit_30.s<3> ;
  assign \sum_4bit_30<2>  = \adder_4bit_30.s<2> ;
  assign \sum_4bit_30<1>  = \adder_4bit_30.s<1> ;
  assign \sum_4bit_30<0>  = \adder_4bit_30.s<0> ;
  assign \sum_4bit_29<4>  = \adder_4bit_29.s<4> ;
  assign \sum_4bit_29<3>  = \adder_4bit_29.s<3> ;
  assign \sum_4bit_29<2>  = \adder_4bit_29.s<2> ;
  assign \sum_4bit_29<1>  = \adder_4bit_29.s<1> ;
  assign \sum_4bit_29<0>  = \adder_4bit_29.s<0> ;
  assign \sum_4bit_28<4>  = \adder_4bit_28.s<4> ;
  assign \sum_4bit_28<3>  = \adder_4bit_28.s<3> ;
  assign \sum_4bit_28<2>  = \adder_4bit_28.s<2> ;
  assign \sum_4bit_28<1>  = \adder_4bit_28.s<1> ;
  assign \sum_4bit_28<0>  = \adder_4bit_28.s<0> ;
  assign \sum_4bit_27<4>  = \adder_4bit_27.s<4> ;
  assign \sum_4bit_27<3>  = \adder_4bit_27.s<3> ;
  assign \sum_4bit_27<2>  = \adder_4bit_27.s<2> ;
  assign \sum_4bit_27<1>  = \adder_4bit_27.s<1> ;
  assign \sum_4bit_27<0>  = \adder_4bit_27.s<0> ;
  assign \sum_4bit_26<4>  = \adder_4bit_26.s<4> ;
  assign \sum_4bit_26<3>  = \adder_4bit_26.s<3> ;
  assign \sum_4bit_26<2>  = \adder_4bit_26.s<2> ;
  assign \sum_4bit_26<1>  = \adder_4bit_26.s<1> ;
  assign \sum_4bit_26<0>  = \adder_4bit_26.s<0> ;
  assign \sum_4bit_25<4>  = \adder_4bit_25.s<4> ;
  assign \sum_4bit_25<3>  = \adder_4bit_25.s<3> ;
  assign \sum_4bit_25<2>  = \adder_4bit_25.s<2> ;
  assign \sum_4bit_25<1>  = \adder_4bit_25.s<1> ;
  assign \sum_4bit_25<0>  = \adder_4bit_25.s<0> ;
  assign \sum_4bit_24<4>  = \adder_4bit_24.s<4> ;
  assign \sum_4bit_24<3>  = \adder_4bit_24.s<3> ;
  assign \sum_4bit_24<2>  = \adder_4bit_24.s<2> ;
  assign \sum_4bit_24<1>  = \adder_4bit_24.s<1> ;
  assign \sum_4bit_24<0>  = \adder_4bit_24.s<0> ;
  assign \sum_4bit_23<4>  = \adder_4bit_23.s<4> ;
  assign \sum_4bit_23<3>  = \adder_4bit_23.s<3> ;
  assign \sum_4bit_23<2>  = \adder_4bit_23.s<2> ;
  assign \sum_4bit_23<1>  = \adder_4bit_23.s<1> ;
  assign \sum_4bit_23<0>  = \adder_4bit_23.s<0> ;
  assign \sum_4bit_22<4>  = \adder_4bit_22.s<4> ;
  assign \sum_4bit_22<3>  = \adder_4bit_22.s<3> ;
  assign \sum_4bit_22<2>  = \adder_4bit_22.s<2> ;
  assign \sum_4bit_22<1>  = \adder_4bit_22.s<1> ;
  assign \sum_4bit_22<0>  = \adder_4bit_22.s<0> ;
  assign \sum_4bit_21<4>  = \adder_4bit_21.s<4> ;
  assign \sum_4bit_21<3>  = \adder_4bit_21.s<3> ;
  assign \sum_4bit_21<2>  = \adder_4bit_21.s<2> ;
  assign \sum_4bit_21<1>  = \adder_4bit_21.s<1> ;
  assign \sum_4bit_21<0>  = \adder_4bit_21.s<0> ;
  assign \sum_4bit_20<4>  = \adder_4bit_20.s<4> ;
  assign \sum_4bit_20<3>  = \adder_4bit_20.s<3> ;
  assign \sum_4bit_20<2>  = \adder_4bit_20.s<2> ;
  assign \sum_4bit_20<1>  = \adder_4bit_20.s<1> ;
  assign \sum_4bit_20<0>  = \adder_4bit_20.s<0> ;
  assign \sum_4bit_19<4>  = \adder_4bit_19.s<4> ;
  assign \sum_4bit_19<3>  = \adder_4bit_19.s<3> ;
  assign \sum_4bit_19<2>  = \adder_4bit_19.s<2> ;
  assign \sum_4bit_19<1>  = \adder_4bit_19.s<1> ;
  assign \sum_4bit_19<0>  = \adder_4bit_19.s<0> ;
  assign \sum_4bit_18<4>  = \adder_4bit_18.s<4> ;
  assign \sum_4bit_18<3>  = \adder_4bit_18.s<3> ;
  assign \sum_4bit_18<2>  = \adder_4bit_18.s<2> ;
  assign \sum_4bit_18<1>  = \adder_4bit_18.s<1> ;
  assign \sum_4bit_18<0>  = \adder_4bit_18.s<0> ;
  assign \sum_4bit_17<4>  = \adder_4bit_17.s<4> ;
  assign \sum_4bit_17<3>  = \adder_4bit_17.s<3> ;
  assign \sum_4bit_17<2>  = \adder_4bit_17.s<2> ;
  assign \sum_4bit_17<1>  = \adder_4bit_17.s<1> ;
  assign \sum_4bit_17<0>  = \adder_4bit_17.s<0> ;
  assign \sum_4bit_16<4>  = \adder_4bit_16.s<4> ;
  assign \sum_4bit_16<3>  = \adder_4bit_16.s<3> ;
  assign \sum_4bit_16<2>  = \adder_4bit_16.s<2> ;
  assign \sum_4bit_16<1>  = \adder_4bit_16.s<1> ;
  assign \sum_4bit_16<0>  = \adder_4bit_16.s<0> ;
  assign \sum_4bit_15<4>  = \adder_4bit_15.s<4> ;
  assign \sum_4bit_15<3>  = \adder_4bit_15.s<3> ;
  assign \sum_4bit_15<2>  = \adder_4bit_15.s<2> ;
  assign \sum_4bit_15<1>  = \adder_4bit_15.s<1> ;
  assign \sum_4bit_15<0>  = \adder_4bit_15.s<0> ;
  assign \sum_4bit_14<4>  = \adder_4bit_14.s<4> ;
  assign \sum_4bit_14<3>  = \adder_4bit_14.s<3> ;
  assign \sum_4bit_14<2>  = \adder_4bit_14.s<2> ;
  assign \sum_4bit_14<1>  = \adder_4bit_14.s<1> ;
  assign \sum_4bit_14<0>  = \adder_4bit_14.s<0> ;
  assign \sum_4bit_13<4>  = \adder_4bit_13.s<4> ;
  assign \sum_4bit_13<3>  = \adder_4bit_13.s<3> ;
  assign \sum_4bit_13<2>  = \adder_4bit_13.s<2> ;
  assign \sum_4bit_13<1>  = \adder_4bit_13.s<1> ;
  assign \sum_4bit_13<0>  = \adder_4bit_13.s<0> ;
  assign \sum_4bit_12<4>  = \adder_4bit_12.s<4> ;
  assign \sum_4bit_12<3>  = \adder_4bit_12.s<3> ;
  assign \sum_4bit_12<2>  = \adder_4bit_12.s<2> ;
  assign \sum_4bit_12<1>  = \adder_4bit_12.s<1> ;
  assign \sum_4bit_12<0>  = \adder_4bit_12.s<0> ;
  assign \sum_4bit_11<4>  = \adder_4bit_11.s<4> ;
  assign \sum_4bit_11<3>  = \adder_4bit_11.s<3> ;
  assign \sum_4bit_11<2>  = \adder_4bit_11.s<2> ;
  assign \sum_4bit_11<1>  = \adder_4bit_11.s<1> ;
  assign \sum_4bit_11<0>  = \adder_4bit_11.s<0> ;
  assign \sum_4bit_10<4>  = \adder_4bit_10.s<4> ;
  assign \sum_4bit_10<3>  = \adder_4bit_10.s<3> ;
  assign \sum_4bit_10<2>  = \adder_4bit_10.s<2> ;
  assign \sum_4bit_10<1>  = \adder_4bit_10.s<1> ;
  assign \sum_4bit_10<0>  = \adder_4bit_10.s<0> ;
  assign \sum_4bit_9<4>  = \adder_4bit_9.s<4> ;
  assign \sum_4bit_9<3>  = \adder_4bit_9.s<3> ;
  assign \sum_4bit_9<2>  = \adder_4bit_9.s<2> ;
  assign \sum_4bit_9<1>  = \adder_4bit_9.s<1> ;
  assign \sum_4bit_9<0>  = \adder_4bit_9.s<0> ;
  assign \sum_4bit_8<4>  = \adder_4bit_8.s<4> ;
  assign \sum_4bit_8<3>  = \adder_4bit_8.s<3> ;
  assign \sum_4bit_8<2>  = \adder_4bit_8.s<2> ;
  assign \sum_4bit_8<1>  = \adder_4bit_8.s<1> ;
  assign \sum_4bit_8<0>  = \adder_4bit_8.s<0> ;
  assign \sum_4bit_7<4>  = \adder_4bit_7.s<4> ;
  assign \sum_4bit_7<3>  = \adder_4bit_7.s<3> ;
  assign \sum_4bit_7<2>  = \adder_4bit_7.s<2> ;
  assign \sum_4bit_7<1>  = \adder_4bit_7.s<1> ;
  assign \sum_4bit_7<0>  = \adder_4bit_7.s<0> ;
  assign \sum_4bit_6<4>  = \adder_4bit_6.s<4> ;
  assign \sum_4bit_6<3>  = \adder_4bit_6.s<3> ;
  assign \sum_4bit_6<2>  = \adder_4bit_6.s<2> ;
  assign \sum_4bit_6<1>  = \adder_4bit_6.s<1> ;
  assign \sum_4bit_6<0>  = \adder_4bit_6.s<0> ;
  assign \sum_4bit_5<4>  = \adder_4bit_5.s<4> ;
  assign \sum_4bit_5<3>  = \adder_4bit_5.s<3> ;
  assign \sum_4bit_5<2>  = \adder_4bit_5.s<2> ;
  assign \sum_4bit_5<1>  = \adder_4bit_5.s<1> ;
  assign \sum_4bit_5<0>  = \adder_4bit_5.s<0> ;
  assign \sum_4bit_4<4>  = \adder_4bit_4.s<4> ;
  assign \sum_4bit_4<3>  = \adder_4bit_4.s<3> ;
  assign \sum_4bit_4<2>  = \adder_4bit_4.s<2> ;
  assign \sum_4bit_4<1>  = \adder_4bit_4.s<1> ;
  assign \sum_4bit_4<0>  = \adder_4bit_4.s<0> ;
  assign \sum_4bit_3<4>  = \adder_4bit_3.s<4> ;
  assign \sum_4bit_3<3>  = \adder_4bit_3.s<3> ;
  assign \sum_4bit_3<2>  = \adder_4bit_3.s<2> ;
  assign \sum_4bit_3<1>  = \adder_4bit_3.s<1> ;
  assign \sum_4bit_3<0>  = \adder_4bit_3.s<0> ;
  assign \sum_4bit_2<4>  = \adder_4bit_2.s<4> ;
  assign \sum_4bit_2<3>  = \adder_4bit_2.s<3> ;
  assign \sum_4bit_2<2>  = \adder_4bit_2.s<2> ;
  assign \sum_4bit_2<1>  = \adder_4bit_2.s<1> ;
  assign \sum_4bit_2<0>  = \adder_4bit_2.s<0> ;
  assign \sum_4bit_1<4>  = \adder_4bit_1.s<4> ;
  assign \sum_4bit_1<3>  = \adder_4bit_1.s<3> ;
  assign \sum_4bit_1<2>  = \adder_4bit_1.s<2> ;
  assign \sum_4bit_1<1>  = \adder_4bit_1.s<1> ;
  assign \sum_4bit_1<0>  = \adder_4bit_1.s<0> ;
  assign \sum_4bit_0<4>  = \adder_4bit_0.s<4> ;
  assign \sum_4bit_0<3>  = \adder_4bit_0.s<3> ;
  assign \sum_4bit_0<2>  = \adder_4bit_0.s<2> ;
  assign \sum_4bit_0<1>  = \adder_4bit_0.s<1> ;
  assign \sum_4bit_0<0>  = \adder_4bit_0.s<0> ;
  assign \out<9>  = \adder_9bit.s<9> ;
  assign \out<8>  = \adder_9bit.s<8> ;
  assign \out<7>  = \adder_9bit.s<7> ;
  assign \out<6>  = \adder_9bit.s<6> ;
  assign \out<5>  = \adder_9bit.s<5> ;
  assign \out<4>  = \adder_9bit.s<4> ;
  assign \out<3>  = \adder_9bit.s<3> ;
  assign \out<2>  = \adder_9bit.s<2> ;
  assign \out<1>  = \adder_9bit.s<1> ;
  assign \out<0>  = \adder_9bit.s<0> ;
  assign \adder_4bit_1.a<3>  = \in_2<3> ;
  assign \adder_4bit_1.a<2>  = \in_2<2> ;
  assign \adder_4bit_1.a<1>  = \in_2<1> ;
  assign \adder_4bit_1.a<0>  = \in_2<0> ;
  assign \adder_4bit_11.b<3>  = \in_23<3> ;
  assign \adder_4bit_11.b<2>  = \in_23<2> ;
  assign \adder_4bit_11.b<1>  = \in_23<1> ;
  assign \adder_4bit_11.b<0>  = \in_23<0> ;
  assign \adder_5bit_7.b<4>  = \adder_4bit_15.s<4> ;
  assign \adder_5bit_7.b<3>  = \adder_4bit_15.s<3> ;
  assign \adder_5bit_7.b<2>  = \adder_4bit_15.s<2> ;
  assign \adder_5bit_7.b<1>  = \adder_4bit_15.s<1> ;
  assign \adder_5bit_7.b<0>  = \adder_4bit_15.s<0> ;
  assign \adder_5bit_6.a<4>  = \adder_4bit_12.s<4> ;
  assign \adder_5bit_6.a<3>  = \adder_4bit_12.s<3> ;
  assign \adder_5bit_6.a<2>  = \adder_4bit_12.s<2> ;
  assign \adder_5bit_6.a<1>  = \adder_4bit_12.s<1> ;
  assign \adder_5bit_6.a<0>  = \adder_4bit_12.s<0> ;
  assign \adder_5bit_6.b<4>  = \adder_4bit_13.s<4> ;
  assign \adder_5bit_6.b<3>  = \adder_4bit_13.s<3> ;
  assign \adder_5bit_6.b<2>  = \adder_4bit_13.s<2> ;
  assign \adder_5bit_6.b<1>  = \adder_4bit_13.s<1> ;
  assign \adder_5bit_6.b<0>  = \adder_4bit_13.s<0> ;
  assign \adder_4bit_20.b<3>  = \in_41<3> ;
  assign \adder_4bit_20.b<2>  = \in_41<2> ;
  assign \adder_4bit_20.b<1>  = \in_41<1> ;
  assign \adder_4bit_20.b<0>  = \in_41<0> ;
  assign \adder_4bit_0.b<3>  = \in_1<3> ;
  assign \adder_4bit_0.b<2>  = \in_1<2> ;
  assign \adder_4bit_0.b<1>  = \in_1<1> ;
  assign \adder_4bit_0.b<0>  = \in_1<0> ;
  assign \adder_5bit_15.a<4>  = \adder_4bit_30.s<4> ;
  assign \adder_5bit_15.a<3>  = \adder_4bit_30.s<3> ;
  assign \adder_5bit_15.a<2>  = \adder_4bit_30.s<2> ;
  assign \adder_5bit_15.a<1>  = \adder_4bit_30.s<1> ;
  assign \adder_5bit_15.a<0>  = \adder_4bit_30.s<0> ;
  assign \adder_5bit_15.b<4>  = \adder_4bit_31.s<4> ;
  assign \adder_5bit_15.b<3>  = \adder_4bit_31.s<3> ;
  assign \adder_5bit_15.b<2>  = \adder_4bit_31.s<2> ;
  assign \adder_5bit_15.b<1>  = \adder_4bit_31.s<1> ;
  assign \adder_5bit_15.b<0>  = \adder_4bit_31.s<0> ;
  assign \adder_5bit_14.a<4>  = \adder_4bit_28.s<4> ;
  assign \adder_5bit_14.a<3>  = \adder_4bit_28.s<3> ;
  assign \adder_5bit_14.a<2>  = \adder_4bit_28.s<2> ;
  assign \adder_5bit_14.a<1>  = \adder_4bit_28.s<1> ;
  assign \adder_5bit_14.a<0>  = \adder_4bit_28.s<0> ;
  assign \adder_5bit_14.b<4>  = \adder_4bit_29.s<4> ;
  assign \adder_5bit_14.b<3>  = \adder_4bit_29.s<3> ;
  assign \adder_5bit_14.b<2>  = \adder_4bit_29.s<2> ;
  assign \adder_5bit_14.b<1>  = \adder_4bit_29.s<1> ;
  assign \adder_5bit_14.b<0>  = \adder_4bit_29.s<0> ;
  assign \adder_4bit_12.a<3>  = \in_24<3> ;
  assign \adder_4bit_12.a<2>  = \in_24<2> ;
  assign \adder_4bit_12.a<1>  = \in_24<1> ;
  assign \adder_4bit_12.a<0>  = \in_24<0> ;
  assign \adder_4bit_12.b<3>  = \in_25<3> ;
  assign \adder_4bit_12.b<2>  = \in_25<2> ;
  assign \adder_4bit_12.b<1>  = \in_25<1> ;
  assign \adder_4bit_12.b<0>  = \in_25<0> ;
  assign \adder_4bit_10.b<3>  = \in_21<3> ;
  assign \adder_4bit_10.b<2>  = \in_21<2> ;
  assign \adder_4bit_10.b<1>  = \in_21<1> ;
  assign \adder_4bit_10.b<0>  = \in_21<0> ;
  assign \adder_5bit_9.b<4>  = \adder_4bit_19.s<4> ;
  assign \adder_5bit_9.b<3>  = \adder_4bit_19.s<3> ;
  assign \adder_5bit_9.b<2>  = \adder_4bit_19.s<2> ;
  assign \adder_5bit_9.b<1>  = \adder_4bit_19.s<1> ;
  assign \adder_5bit_9.b<0>  = \adder_4bit_19.s<0> ;
  assign \adder_5bit_8.b<4>  = \adder_4bit_17.s<4> ;
  assign \adder_5bit_8.b<3>  = \adder_4bit_17.s<3> ;
  assign \adder_5bit_8.b<2>  = \adder_4bit_17.s<2> ;
  assign \adder_5bit_8.b<1>  = \adder_4bit_17.s<1> ;
  assign \adder_5bit_8.b<0>  = \adder_4bit_17.s<0> ;
  assign \adder_4bit_14.a<3>  = \in_28<3> ;
  assign \adder_4bit_14.a<2>  = \in_28<2> ;
  assign \adder_4bit_14.a<1>  = \in_28<1> ;
  assign \adder_4bit_14.a<0>  = \in_28<0> ;
  assign \adder_4bit_14.b<3>  = \in_29<3> ;
  assign \adder_4bit_14.b<2>  = \in_29<2> ;
  assign \adder_4bit_14.b<1>  = \in_29<1> ;
  assign \adder_4bit_14.b<0>  = \in_29<0> ;
  assign \adder_4bit_21.b<3>  = \in_43<3> ;
  assign \adder_4bit_21.b<2>  = \in_43<2> ;
  assign \adder_4bit_21.b<1>  = \in_43<1> ;
  assign \adder_4bit_21.b<0>  = \in_43<0> ;
  assign \adder_4bit_31.a<3>  = \in_62<3> ;
  assign \adder_4bit_31.a<2>  = \in_62<2> ;
  assign \adder_4bit_31.a<1>  = \in_62<1> ;
  assign \adder_4bit_31.a<0>  = \in_62<0> ;
  assign \adder_4bit_31.b<3>  = \in_63<3> ;
  assign \adder_4bit_31.b<2>  = \in_63<2> ;
  assign \adder_4bit_31.b<1>  = \in_63<1> ;
  assign \adder_4bit_31.b<0>  = \in_63<0> ;
  assign \adder_4bit_25.b<3>  = \in_51<3> ;
  assign \adder_4bit_25.b<2>  = \in_51<2> ;
  assign \adder_4bit_25.b<1>  = \in_51<1> ;
  assign \adder_4bit_25.b<0>  = \in_51<0> ;
  assign \adder_4bit_9.b<3>  = \in_19<3> ;
  assign \adder_4bit_9.b<2>  = \in_19<2> ;
  assign \adder_4bit_9.b<1>  = \in_19<1> ;
  assign \adder_4bit_9.b<0>  = \in_19<0> ;
  assign \adder_5bit_11.b<4>  = \adder_4bit_23.s<4> ;
  assign \adder_5bit_11.b<3>  = \adder_4bit_23.s<3> ;
  assign \adder_5bit_11.b<2>  = \adder_4bit_23.s<2> ;
  assign \adder_5bit_11.b<1>  = \adder_4bit_23.s<1> ;
  assign \adder_5bit_11.b<0>  = \adder_4bit_23.s<0> ;
  assign \adder_5bit_10.b<4>  = \adder_4bit_21.s<4> ;
  assign \adder_5bit_10.b<3>  = \adder_4bit_21.s<3> ;
  assign \adder_5bit_10.b<2>  = \adder_4bit_21.s<2> ;
  assign \adder_5bit_10.b<1>  = \adder_4bit_21.s<1> ;
  assign \adder_5bit_10.b<0>  = \adder_4bit_21.s<0> ;
  assign \adder_4bit_26.b<3>  = \in_53<3> ;
  assign \adder_4bit_26.b<2>  = \in_53<2> ;
  assign \adder_4bit_26.b<1>  = \in_53<1> ;
  assign \adder_4bit_26.b<0>  = \in_53<0> ;
  assign \adder_4bit_24.a<3>  = \in_48<3> ;
  assign \adder_4bit_24.a<2>  = \in_48<2> ;
  assign \adder_4bit_24.a<1>  = \in_48<1> ;
  assign \adder_4bit_24.a<0>  = \in_48<0> ;
  assign \adder_4bit_24.b<3>  = \in_49<3> ;
  assign \adder_4bit_24.b<2>  = \in_49<2> ;
  assign \adder_4bit_24.b<1>  = \in_49<1> ;
  assign \adder_4bit_24.b<0>  = \in_49<0> ;
  assign \adder_4bit_28.a<3>  = \in_56<3> ;
  assign \adder_4bit_28.a<2>  = \in_56<2> ;
  assign \adder_4bit_28.a<1>  = \in_56<1> ;
  assign \adder_4bit_28.a<0>  = \in_56<0> ;
  assign \adder_4bit_28.b<3>  = \in_57<3> ;
  assign \adder_4bit_28.b<2>  = \in_57<2> ;
  assign \adder_4bit_28.b<1>  = \in_57<1> ;
  assign \adder_4bit_28.b<0>  = \in_57<0> ;
  assign \adder_5bit_3.b<4>  = \adder_4bit_7.s<4> ;
  assign \adder_5bit_3.b<3>  = \adder_4bit_7.s<3> ;
  assign \adder_5bit_3.b<2>  = \adder_4bit_7.s<2> ;
  assign \adder_5bit_3.b<1>  = \adder_4bit_7.s<1> ;
  assign \adder_5bit_3.b<0>  = \adder_4bit_7.s<0> ;
  assign \adder_4bit_1.b<3>  = \in_3<3> ;
  assign \adder_4bit_1.b<2>  = \in_3<2> ;
  assign \adder_4bit_1.b<1>  = \in_3<1> ;
  assign \adder_4bit_1.b<0>  = \in_3<0> ;
  assign \adder_4bit_8.b<3>  = \in_17<3> ;
  assign \adder_4bit_8.b<2>  = \in_17<2> ;
  assign \adder_4bit_8.b<1>  = \in_17<1> ;
  assign \adder_4bit_8.b<0>  = \in_17<0> ;
  assign \adder_4bit_5.a<3>  = \in_10<3> ;
  assign \adder_4bit_5.a<2>  = \in_10<2> ;
  assign \adder_4bit_5.a<1>  = \in_10<1> ;
  assign \adder_4bit_5.a<0>  = \in_10<0> ;
  assign \adder_4bit_0.a<3>  = \in_0<3> ;
  assign \adder_4bit_0.a<2>  = \in_0<2> ;
  assign \adder_4bit_0.a<1>  = \in_0<1> ;
  assign \adder_4bit_0.a<0>  = \in_0<0> ;
  assign \adder_4bit_4.a<3>  = \in_8<3> ;
  assign \adder_4bit_4.a<2>  = \in_8<2> ;
  assign \adder_4bit_4.a<1>  = \in_8<1> ;
  assign \adder_4bit_4.a<0>  = \in_8<0> ;
  assign \adder_4bit_7.a<3>  = \in_14<3> ;
  assign \adder_4bit_7.a<2>  = \in_14<2> ;
  assign \adder_4bit_7.a<1>  = \in_14<1> ;
  assign \adder_4bit_7.a<0>  = \in_14<0> ;
  assign \adder_4bit_7.b<3>  = \in_15<3> ;
  assign \adder_4bit_7.b<2>  = \in_15<2> ;
  assign \adder_4bit_7.b<1>  = \in_15<1> ;
  assign \adder_4bit_7.b<0>  = \in_15<0> ;
  assign \adder_4bit_3.a<3>  = \in_6<3> ;
  assign \adder_4bit_3.a<2>  = \in_6<2> ;
  assign \adder_4bit_3.a<1>  = \in_6<1> ;
  assign \adder_4bit_3.a<0>  = \in_6<0> ;
  assign \adder_9bit.sign  = sign_weight;
  assign \adder_8bit_1.sign  = sign_weight;
  assign \adder_4bit_13.b<3>  = \in_27<3> ;
  assign \adder_4bit_13.b<2>  = \in_27<2> ;
  assign \adder_8bit_0.sign  = sign_weight;
  assign \adder_4bit_13.b<0>  = \in_27<0> ;
  assign \adder_5bit_2.b<4>  = \adder_4bit_5.s<4> ;
  assign \adder_4bit_13.b<1>  = \in_27<1> ;
  assign \adder_7bit_3.sign  = sign_weight;
  assign \adder_5bit_2.b<2>  = \adder_4bit_5.s<2> ;
  assign \adder_5bit_2.b<3>  = \adder_4bit_5.s<3> ;
  assign \adder_5bit_2.b<1>  = \adder_4bit_5.s<1> ;
  assign \adder_7bit_2.sign  = sign_weight;
  assign \adder_5bit_2.b<0>  = \adder_4bit_5.s<0> ;
  assign \adder_7bit_1.sign  = sign_weight;
  assign \adder_7bit_0.sign  = sign_weight;
  assign \adder_4bit_2.a<0>  = \in_4<0> ;
  assign \adder_6bit_7.sign  = sign_weight;
  assign \adder_5bit_5.a<3>  = \adder_4bit_10.s<3> ;
  assign \adder_5bit_5.a<4>  = \adder_4bit_10.s<4> ;
  assign \adder_5bit_5.a<2>  = \adder_4bit_10.s<2> ;
  assign \adder_6bit_6.sign  = sign_weight;
  assign \adder_5bit_5.a<0>  = \adder_4bit_10.s<0> ;
  assign \adder_5bit_5.b<4>  = \adder_4bit_11.s<4> ;
  assign \adder_5bit_5.a<1>  = \adder_4bit_10.s<1> ;
  assign \adder_5bit_5.b<3>  = \adder_4bit_11.s<3> ;
  assign \adder_6bit_5.sign  = sign_weight;
  assign \adder_4bit_16.b<0>  = \in_33<0> ;
  assign \adder_4bit_17.a<3>  = \in_34<3> ;
  assign \adder_5bit_5.b<2>  = \adder_4bit_11.s<2> ;
  assign \adder_5bit_5.b<1>  = \adder_4bit_11.s<1> ;
  assign \adder_6bit_4.sign  = sign_weight;
  assign \adder_5bit_4.a<4>  = \adder_4bit_8.s<4> ;
  assign \adder_5bit_4.a<3>  = \adder_4bit_8.s<3> ;
  assign \adder_5bit_5.b<0>  = \adder_4bit_11.s<0> ;
  assign \adder_5bit_4.a<2>  = \adder_4bit_8.s<2> ;
  assign \adder_6bit_3.sign  = sign_weight;
  assign \adder_5bit_4.a<0>  = \adder_4bit_8.s<0> ;
  assign \adder_5bit_4.b<4>  = \adder_4bit_9.s<4> ;
  assign \adder_5bit_4.a<1>  = \adder_4bit_8.s<1> ;
  assign \adder_5bit_4.b<3>  = \adder_4bit_9.s<3> ;
  assign \adder_6bit_2.sign  = sign_weight;
  assign \adder_5bit_1.b<4>  = \adder_4bit_3.s<4> ;
  assign \adder_5bit_1.b<3>  = \adder_4bit_3.s<3> ;
  assign \adder_5bit_4.b<2>  = \adder_4bit_9.s<2> ;
  assign \adder_5bit_4.b<1>  = \adder_4bit_9.s<1> ;
  assign \adder_6bit_1.sign  = sign_weight;
  assign \adder_5bit_1.b<2>  = \adder_4bit_3.s<2> ;
  assign \adder_5bit_1.b<1>  = \adder_4bit_3.s<1> ;
  assign \adder_5bit_4.b<0>  = \adder_4bit_9.s<0> ;
  assign \adder_6bit_2.a<5>  = \adder_5bit_4.s<5> ;
  assign \adder_6bit_0.sign  = sign_weight;
  assign \adder_6bit_2.a<3>  = \adder_5bit_4.s<3> ;
  assign \adder_5bit_1.b<0>  = \adder_4bit_3.s<0> ;
  assign \adder_6bit_2.a<4>  = \adder_5bit_4.s<4> ;
  assign \adder_6bit_2.a<2>  = \adder_5bit_4.s<2> ;
  assign \adder_5bit_15.sign  = sign_weight;
  assign \adder_6bit_2.a<1>  = \adder_5bit_4.s<1> ;
  assign \adder_6bit_2.b<5>  = \adder_5bit_5.s<5> ;
  assign \adder_5bit_14.sign  = sign_weight;
  assign \adder_6bit_2.a<0>  = \adder_5bit_4.s<0> ;
  assign \adder_6bit_2.b<3>  = \adder_5bit_5.s<3> ;
  assign \adder_5bit_13.sign  = sign_weight;
  assign \adder_6bit_2.b<2>  = \adder_5bit_5.s<2> ;
  assign \adder_4bit_15.b<3>  = \in_31<3> ;
  assign \adder_6bit_2.b<4>  = \adder_5bit_5.s<4> ;
  assign \adder_4bit_15.b<2>  = \in_31<2> ;
  assign \adder_5bit_12.sign  = sign_weight;
  assign \adder_4bit_15.b<1>  = \in_31<1> ;
  assign \adder_4bit_15.b<0>  = \in_31<0> ;
  assign \adder_6bit_2.b<1>  = \adder_5bit_5.s<1> ;
  assign \adder_6bit_1.a<5>  = \adder_5bit_2.s<5> ;
  assign \adder_5bit_11.sign  = sign_weight;
  assign \adder_6bit_1.a<4>  = \adder_5bit_2.s<4> ;
  assign \adder_7bit_2.b<5>  = \adder_6bit_5.s<5> ;
  assign \adder_6bit_2.b<0>  = \adder_5bit_5.s<0> ;
  assign \adder_6bit_1.a<2>  = \adder_5bit_2.s<2> ;
  assign \adder_5bit_10.sign  = sign_weight;
  assign \adder_6bit_1.a<1>  = \adder_5bit_2.s<1> ;
  assign \adder_7bit_2.b<4>  = \adder_6bit_5.s<4> ;
  assign \adder_6bit_1.a<3>  = \adder_5bit_2.s<3> ;
  assign \adder_6bit_1.b<5>  = \adder_5bit_3.s<5> ;
  assign \adder_5bit_9.sign  = sign_weight;
  assign \adder_6bit_1.b<4>  = \adder_5bit_3.s<4> ;
  assign \adder_6bit_1.a<0>  = \adder_5bit_2.s<0> ;
  assign \adder_6bit_1.b<2>  = \adder_5bit_3.s<2> ;
  assign \adder_5bit_8.sign  = sign_weight;
  assign \adder_6bit_1.b<1>  = \adder_5bit_3.s<1> ;
  assign \adder_6bit_1.b<3>  = \adder_5bit_3.s<3> ;
  assign \adder_6bit_0.b<5>  = \adder_5bit_1.s<5> ;
  assign \adder_5bit_7.sign  = sign_weight;
  assign \adder_6bit_0.b<4>  = \adder_5bit_1.s<4> ;
  assign \adder_7bit_3.a<3>  = \adder_6bit_6.s<3> ;
  assign \adder_6bit_1.b<0>  = \adder_5bit_3.s<0> ;
  assign \adder_7bit_3.a<2>  = \adder_6bit_6.s<2> ;
  assign \adder_5bit_6.sign  = sign_weight;
  assign \adder_7bit_3.a<1>  = \adder_6bit_6.s<1> ;
  assign \adder_7bit_3.a<0>  = \adder_6bit_6.s<0> ;
  assign \adder_6bit_0.b<3>  = \adder_5bit_1.s<3> ;
  assign \adder_4bit_2.b<0>  = \in_5<0> ;
  assign \adder_5bit_5.sign  = sign_weight;
  assign \adder_4bit_27.b<3>  = \in_55<3> ;
  assign \adder_4bit_27.b<2>  = \in_55<2> ;
  assign \adder_6bit_0.b<2>  = \adder_5bit_1.s<2> ;
  assign \adder_6bit_0.b<0>  = \adder_5bit_1.s<0> ;
  assign \adder_5bit_4.sign  = sign_weight;
  assign \adder_4bit_27.b<1>  = \in_55<1> ;
  assign \adder_4bit_27.b<0>  = \in_55<0> ;
  assign \adder_6bit_0.b<1>  = \adder_5bit_1.s<1> ;
  assign \adder_5bit_13.b<3>  = \adder_4bit_27.s<3> ;
  assign \adder_5bit_3.sign  = sign_weight;
  assign \adder_5bit_13.b<2>  = \adder_4bit_27.s<2> ;
  assign \adder_5bit_13.b<4>  = \adder_4bit_27.s<4> ;
  assign \adder_5bit_13.b<0>  = \adder_4bit_27.s<0> ;
  assign \adder_5bit_2.sign  = sign_weight;
  assign \adder_4bit_2.b<2>  = \in_5<2> ;
  assign \adder_5bit_13.b<1>  = \adder_4bit_27.s<1> ;
  assign \adder_4bit_2.a<1>  = \in_4<1> ;
  assign \adder_5bit_1.sign  = sign_weight;
  assign \adder_4bit_6.a<1>  = \in_12<1> ;
  assign \adder_4bit_2.b<1>  = \in_5<1> ;
  assign \adder_5bit_0.sign  = sign_weight;
  assign \adder_5bit_12.a<4>  = \adder_4bit_24.s<4> ;
  assign \adder_4bit_31.sign  = sign_weight;
  assign \adder_7bit_2.a<3>  = \adder_6bit_4.s<3> ;
  assign \adder_7bit_2.a<2>  = \adder_6bit_4.s<2> ;
  assign \adder_5bit_12.a<3>  = \adder_4bit_24.s<3> ;
  assign \adder_5bit_12.a<1>  = \adder_4bit_24.s<1> ;
  assign \adder_4bit_30.sign  = sign_weight;
  assign \adder_5bit_12.a<0>  = \adder_4bit_24.s<0> ;
  assign \adder_4bit_17.a<1>  = \in_34<1> ;
  assign \adder_5bit_12.a<2>  = \adder_4bit_24.s<2> ;
  assign \adder_5bit_12.b<3>  = \adder_4bit_25.s<3> ;
  assign \adder_4bit_29.sign  = sign_weight;
  assign \adder_5bit_12.b<2>  = \adder_4bit_25.s<2> ;
  assign \adder_4bit_17.a<0>  = \in_34<0> ;
  assign \adder_5bit_12.b<4>  = \adder_4bit_25.s<4> ;
  assign \adder_4bit_28.sign  = sign_weight;
  assign \adder_5bit_12.b<1>  = \adder_4bit_25.s<1> ;
  assign \adder_4bit_27.sign  = sign_weight;
  assign \adder_5bit_12.b<0>  = \adder_4bit_25.s<0> ;
  assign \adder_4bit_26.sign  = sign_weight;
  assign \adder_4bit_6.a<3>  = \in_12<3> ;
  assign \adder_7bit_2.b<3>  = \adder_6bit_5.s<3> ;
  assign \adder_7bit_2.a<1>  = \adder_6bit_4.s<1> ;
  assign \adder_4bit_25.sign  = sign_weight;
  assign \adder_4bit_6.a<0>  = \in_12<0> ;
  assign \adder_7bit_2.a<0>  = \adder_6bit_4.s<0> ;
  assign \adder_4bit_6.a<2>  = \in_12<2> ;
  assign \adder_4bit_6.b<2>  = \in_13<2> ;
  assign \adder_4bit_24.sign  = sign_weight;
  assign \adder_7bit_2.b<1>  = \adder_6bit_5.s<1> ;
  assign \adder_7bit_2.b<0>  = \adder_6bit_5.s<0> ;
  assign \adder_4bit_6.b<3>  = \in_13<3> ;
  assign \adder_4bit_6.b<0>  = \in_13<0> ;
  assign \adder_4bit_23.sign  = sign_weight;
  assign \adder_6bit_5.a<5>  = \adder_5bit_10.s<5> ;
  assign \adder_4bit_17.a<2>  = \in_34<2> ;
  assign \adder_4bit_6.b<1>  = \in_13<1> ;
  assign \adder_4bit_17.b<3>  = \in_35<3> ;
  assign \adder_4bit_22.sign  = sign_weight;
  assign \adder_4bit_17.b<1>  = \in_35<1> ;
  assign \adder_4bit_17.b<2>  = \in_35<2> ;
  assign \adder_6bit_5.a<4>  = \adder_5bit_10.s<4> ;
  assign \adder_6bit_5.a<2>  = \adder_5bit_10.s<2> ;
  assign \adder_4bit_21.sign  = sign_weight;
  assign \adder_6bit_5.a<1>  = \adder_5bit_10.s<1> ;
  assign \adder_7bit_2.a<5>  = \adder_6bit_4.s<5> ;
  assign \adder_6bit_5.a<3>  = \adder_5bit_10.s<3> ;
  assign \adder_6bit_5.b<5>  = \adder_5bit_11.s<5> ;
  assign \adder_4bit_20.sign  = sign_weight;
  assign \adder_6bit_5.b<4>  = \adder_5bit_11.s<4> ;
  assign \adder_6bit_5.a<0>  = \adder_5bit_10.s<0> ;
  assign \adder_6bit_5.b<2>  = \adder_5bit_11.s<2> ;
  assign \adder_4bit_19.sign  = sign_weight;
  assign \adder_6bit_5.b<1>  = \adder_5bit_11.s<1> ;
  assign \adder_6bit_5.b<3>  = \adder_5bit_11.s<3> ;
  assign \adder_4bit_23.b<2>  = \in_47<2> ;
  assign \adder_4bit_18.sign  = sign_weight;
  assign \adder_6bit_5.b<0>  = \adder_5bit_11.s<0> ;
  assign \adder_4bit_23.b<1>  = \in_47<1> ;
  assign \adder_4bit_17.sign  = sign_weight;
  assign \adder_4bit_2.a<3>  = \in_4<3> ;
  assign \adder_4bit_2.a<2>  = \in_4<2> ;
  assign \adder_4bit_23.b<3>  = \in_47<3> ;
  assign \adder_4bit_30.b<3>  = \in_61<3> ;
  assign \adder_4bit_16.sign  = sign_weight;
  assign \adder_4bit_30.b<2>  = \in_61<2> ;
  assign \adder_4bit_23.b<0>  = \in_47<0> ;
  assign \adder_4bit_30.b<0>  = \in_61<0> ;
  assign \adder_4bit_15.sign  = sign_weight;
  assign \adder_4bit_29.b<3>  = \in_59<3> ;
  assign \adder_4bit_30.b<1>  = \in_61<1> ;
  assign \adder_4bit_29.b<1>  = \in_59<1> ;
  assign \adder_4bit_14.sign  = sign_weight;
  assign \adder_7bit_2.a<6>  = \adder_6bit_4.s<6> ;
  assign \adder_4bit_29.b<2>  = \in_59<2> ;
  assign \adder_4bit_13.sign  = sign_weight;
  assign \adder_4bit_2.b<3>  = \in_5<3> ;
  assign \adder_4bit_29.b<0>  = \in_59<0> ;
  assign \adder_4bit_12.sign  = sign_weight;
  assign \adder_4bit_22.b<3>  = \in_45<3> ;
  assign \adder_4bit_11.sign  = sign_weight;
  assign \adder_4bit_22.b<2>  = \in_45<2> ;
  assign \adder_7bit_3.a<4>  = \adder_6bit_6.s<4> ;
  assign \adder_4bit_22.b<0>  = \in_45<0> ;
  assign \adder_4bit_10.sign  = sign_weight;
  assign \adder_4bit_22.a<3>  = \in_44<3> ;
  assign \adder_4bit_22.b<1>  = \in_45<1> ;
  assign \adder_4bit_22.a<1>  = \in_44<1> ;
  assign \adder_4bit_9.sign  = sign_weight;
  assign \adder_4bit_22.a<0>  = \in_44<0> ;
  assign \adder_7bit_2.b<6>  = \adder_6bit_5.s<6> ;
  assign \adder_4bit_22.a<2>  = \in_44<2> ;
  assign \adder_4bit_8.sign  = sign_weight;
  assign \adder_4bit_7.sign  = sign_weight;
  assign \adder_4bit_16.b<3>  = \in_33<3> ;
  assign \adder_4bit_6.sign  = sign_weight;
  assign \adder_4bit_16.b<2>  = \in_33<2> ;
  assign \adder_4bit_16.b<1>  = \in_33<1> ;
  assign \adder_4bit_5.b<3>  = \in_11<3> ;
  assign \adder_4bit_17.b<0>  = \in_35<0> ;
  assign \adder_4bit_5.sign  = sign_weight;
  assign \adder_4bit_5.b<2>  = \in_11<2> ;
  assign \adder_4bit_5.b<0>  = \in_11<0> ;
  assign \adder_4bit_4.sign  = sign_weight;
  assign \adder_4bit_5.b<1>  = \in_11<1> ;
  assign \adder_7bit_2.b<2>  = \adder_6bit_5.s<2> ;
  assign \adder_4bit_3.sign  = sign_weight;
  assign \adder_4bit_3.b<3>  = \in_7<3> ;
  assign \adder_4bit_4.b<3>  = \in_9<3> ;
  assign \adder_4bit_3.b<2>  = \in_7<2> ;
  assign \adder_4bit_2.sign  = sign_weight;
  assign \adder_4bit_3.b<1>  = \in_7<1> ;
  assign \adder_4bit_3.b<0>  = \in_7<0> ;
  assign \adder_4bit_4.b<2>  = \in_9<2> ;
  assign \adder_4bit_1.sign  = sign_weight;
  assign \adder_4bit_4.b<1>  = \in_9<1> ;
  assign \adder_4bit_0.sign  = sign_weight;
  assign \adder_7bit_2.a<4>  = \adder_6bit_4.s<4> ;
  assign \adder_4bit_4.b<0>  = \in_9<0> ;
  assign \adder_4bit_18.a<3>  = \in_36<3> ;
  assign \adder_4bit_18.a<2>  = \in_36<2> ;
  assign \adder_4bit_18.a<1>  = \in_36<1> ;
  assign \adder_4bit_18.a<0>  = \in_36<0> ;
  assign \adder_4bit_18.b<3>  = \in_37<3> ;
  assign \adder_4bit_18.b<2>  = \in_37<2> ;
  assign \adder_4bit_18.b<1>  = \in_37<1> ;
  assign \adder_4bit_18.b<0>  = \in_37<0> ;
  assign \adder_4bit_19.b<3>  = \in_39<3> ;
  assign \adder_4bit_19.b<2>  = \in_39<2> ;
  assign \adder_4bit_19.b<1>  = \in_39<1> ;
  assign \adder_4bit_19.b<0>  = \in_39<0> ;
  assign \adder_6bit_7.b<5>  = \adder_5bit_15.s<5> ;
  assign \adder_6bit_7.b<4>  = \adder_5bit_15.s<4> ;
  assign \adder_6bit_7.b<3>  = \adder_5bit_15.s<3> ;
  assign \adder_6bit_7.b<2>  = \adder_5bit_15.s<2> ;
  assign \adder_6bit_7.b<1>  = \adder_5bit_15.s<1> ;
  assign \adder_6bit_7.b<0>  = \adder_5bit_15.s<0> ;
  assign \adder_7bit_3.b<6>  = \adder_6bit_7.s<6> ;
  assign \adder_7bit_3.b<5>  = \adder_6bit_7.s<5> ;
  assign \adder_7bit_3.b<4>  = \adder_6bit_7.s<4> ;
  assign \adder_7bit_3.b<3>  = \adder_6bit_7.s<3> ;
  assign \adder_7bit_3.b<2>  = \adder_6bit_7.s<2> ;
  assign \adder_7bit_3.b<1>  = \adder_6bit_7.s<1> ;
  assign \adder_7bit_3.b<0>  = \adder_6bit_7.s<0> ;
  assign \adder_9bit.a<8>  = \adder_8bit_0.s<8> ;
  assign \adder_9bit.a<7>  = \adder_8bit_0.s<7> ;
  assign \adder_9bit.a<6>  = \adder_8bit_0.s<6> ;
  assign \adder_9bit.a<5>  = \adder_8bit_0.s<5> ;
  assign \adder_9bit.a<4>  = \adder_8bit_0.s<4> ;
  assign \adder_9bit.a<3>  = \adder_8bit_0.s<3> ;
  assign \adder_9bit.a<2>  = \adder_8bit_0.s<2> ;
  assign \adder_9bit.a<1>  = \adder_8bit_0.s<1> ;
  assign \adder_9bit.a<0>  = \adder_8bit_0.s<0> ;
  assign \adder_9bit.b<8>  = \adder_8bit_1.s<8> ;
  assign \adder_9bit.b<7>  = \adder_8bit_1.s<7> ;
  assign \adder_9bit.b<6>  = \adder_8bit_1.s<6> ;
  assign \adder_9bit.b<5>  = \adder_8bit_1.s<5> ;
  assign \adder_9bit.b<4>  = \adder_8bit_1.s<4> ;
  assign \adder_9bit.b<3>  = \adder_8bit_1.s<3> ;
  assign \adder_9bit.b<2>  = \adder_8bit_1.s<2> ;
  assign \adder_9bit.b<1>  = \adder_8bit_1.s<1> ;
  assign \adder_9bit.b<0>  = \adder_8bit_1.s<0> ;
  assign \adder_8bit_1.a<7>  = \adder_7bit_2.s<7> ;
  assign \adder_8bit_1.a<6>  = \adder_7bit_2.s<6> ;
  assign \adder_8bit_1.a<5>  = \adder_7bit_2.s<5> ;
  assign \adder_8bit_1.a<4>  = \adder_7bit_2.s<4> ;
  assign \adder_8bit_1.a<3>  = \adder_7bit_2.s<3> ;
  assign \adder_8bit_1.a<2>  = \adder_7bit_2.s<2> ;
  assign \adder_8bit_1.a<1>  = \adder_7bit_2.s<1> ;
  assign \adder_8bit_1.a<0>  = \adder_7bit_2.s<0> ;
  assign \adder_8bit_1.b<7>  = \adder_7bit_3.s<7> ;
  assign \adder_8bit_1.b<6>  = \adder_7bit_3.s<6> ;
  assign \adder_8bit_1.b<5>  = \adder_7bit_3.s<5> ;
  assign \adder_8bit_1.b<4>  = \adder_7bit_3.s<4> ;
  assign \adder_8bit_1.b<3>  = \adder_7bit_3.s<3> ;
  assign \adder_8bit_1.b<2>  = \adder_7bit_3.s<2> ;
  assign \adder_8bit_1.b<1>  = \adder_7bit_3.s<1> ;
  assign \adder_8bit_1.b<0>  = \adder_7bit_3.s<0> ;
  assign \adder_8bit_0.a<3>  = \adder_7bit_0.s<3> ;
  assign \adder_8bit_0.a<2>  = \adder_7bit_0.s<2> ;
  assign \adder_8bit_0.a<4>  = \adder_7bit_0.s<4> ;
  assign \adder_8bit_0.a<1>  = \adder_7bit_0.s<1> ;
  assign \adder_8bit_0.a<0>  = \adder_7bit_0.s<0> ;
  assign \adder_8bit_0.b<7>  = \adder_7bit_1.s<7> ;
  assign \adder_8bit_0.b<6>  = \adder_7bit_1.s<6> ;
  assign \adder_8bit_0.b<5>  = \adder_7bit_1.s<5> ;
  assign \adder_8bit_0.b<4>  = \adder_7bit_1.s<4> ;
  assign \adder_8bit_0.b<3>  = \adder_7bit_1.s<3> ;
  assign \adder_8bit_0.b<2>  = \adder_7bit_1.s<2> ;
  assign \adder_8bit_0.b<1>  = \adder_7bit_1.s<1> ;
  assign \adder_8bit_0.b<0>  = \adder_7bit_1.s<0> ;
  assign \adder_7bit_3.a<6>  = \adder_6bit_6.s<6> ;
  assign \adder_7bit_3.a<5>  = \adder_6bit_6.s<5> ;
  assign \adder_8bit_0.a<7>  = \adder_7bit_0.s<7> ;
  assign \adder_8bit_0.a<6>  = \adder_7bit_0.s<6> ;
  assign \adder_8bit_0.a<5>  = \adder_7bit_0.s<5> ;
endmodule
