
module decoder_6_to_64(enable, \in<0> , \in<1> , \in<2> , \in<3> , \in<4> , \in<5> , \out<0> , \out<1> , \out<2> , \out<3> , \out<4> , \out<5> , \out<6> , \out<7> , \out<8> , \out<9> , \out<10> , \out<11> , \out<12> , \out<13> , \out<14> , \out<15> , \out<16> , \out<17> , \out<18> , \out<19> , \out<20> , \out<21> , \out<22> , \out<23> , \out<24> , \out<25> , \out<26> , \out<27> , \out<28> , \out<29> , \out<30> , \out<31> , \out<32> , \out<33> , \out<34> , \out<35> , \out<36> , \out<37> , \out<38> , \out<39> , \out<40> , \out<41> , \out<42> , \out<43> , \out<44> , \out<45> , \out<46> , \out<47> , \out<48> , \out<49> , \out<50> , \out<51> , \out<52> , \out<53> , \out<54> , \out<55> , \out<56> , \out<57> , \out<58> , \out<59> , \out<60> , \out<61> , \out<62> , \out<63> );
  input enable;
  input \in<0> ;
  input \in<1> ;
  input \in<2> ;
  input \in<3> ;
  input \in<4> ;
  input \in<5> ;
  wire \in_b<0> ;
  wire \in_b<1> ;
  wire \in_b<2> ;
  wire \in_b<3> ;
  wire \in_b<4> ;
  wire \in_b<5> ;
  wire \nand_0.and_0 ;
  wire \nand_0.and_1 ;
  wire \nand_0.and_2 ;
  wire \nand_0.and_3 ;
  wire \nand_0.and_4 ;
  wire \nand_0.in_0 ;
  wire \nand_0.in_1 ;
  wire \nand_0.in_2 ;
  wire \nand_0.in_3 ;
  wire \nand_0.in_4 ;
  wire \nand_0.in_5 ;
  wire \nand_0.in_6 ;
  wire \nand_0.nand_0 ;
  wire \nand_0.nand_1 ;
  wire \nand_0.nand_2 ;
  wire \nand_0.nand_3 ;
  wire \nand_0.nand_4 ;
  wire \nand_0.out ;
  wire \nand_1.and_0 ;
  wire \nand_1.and_1 ;
  wire \nand_1.and_2 ;
  wire \nand_1.and_3 ;
  wire \nand_1.and_4 ;
  wire \nand_1.in_0 ;
  wire \nand_1.in_1 ;
  wire \nand_1.in_2 ;
  wire \nand_1.in_3 ;
  wire \nand_1.in_4 ;
  wire \nand_1.in_5 ;
  wire \nand_1.in_6 ;
  wire \nand_1.nand_0 ;
  wire \nand_1.nand_1 ;
  wire \nand_1.nand_2 ;
  wire \nand_1.nand_3 ;
  wire \nand_1.nand_4 ;
  wire \nand_1.out ;
  wire \nand_10.and_0 ;
  wire \nand_10.and_1 ;
  wire \nand_10.and_2 ;
  wire \nand_10.and_3 ;
  wire \nand_10.and_4 ;
  wire \nand_10.in_0 ;
  wire \nand_10.in_1 ;
  wire \nand_10.in_2 ;
  wire \nand_10.in_3 ;
  wire \nand_10.in_4 ;
  wire \nand_10.in_5 ;
  wire \nand_10.in_6 ;
  wire \nand_10.nand_0 ;
  wire \nand_10.nand_1 ;
  wire \nand_10.nand_2 ;
  wire \nand_10.nand_3 ;
  wire \nand_10.nand_4 ;
  wire \nand_10.out ;
  wire \nand_11.and_0 ;
  wire \nand_11.and_1 ;
  wire \nand_11.and_2 ;
  wire \nand_11.and_3 ;
  wire \nand_11.and_4 ;
  wire \nand_11.in_0 ;
  wire \nand_11.in_1 ;
  wire \nand_11.in_2 ;
  wire \nand_11.in_3 ;
  wire \nand_11.in_4 ;
  wire \nand_11.in_5 ;
  wire \nand_11.in_6 ;
  wire \nand_11.nand_0 ;
  wire \nand_11.nand_1 ;
  wire \nand_11.nand_2 ;
  wire \nand_11.nand_3 ;
  wire \nand_11.nand_4 ;
  wire \nand_11.out ;
  wire \nand_12.and_0 ;
  wire \nand_12.and_1 ;
  wire \nand_12.and_2 ;
  wire \nand_12.and_3 ;
  wire \nand_12.and_4 ;
  wire \nand_12.in_0 ;
  wire \nand_12.in_1 ;
  wire \nand_12.in_2 ;
  wire \nand_12.in_3 ;
  wire \nand_12.in_4 ;
  wire \nand_12.in_5 ;
  wire \nand_12.in_6 ;
  wire \nand_12.nand_0 ;
  wire \nand_12.nand_1 ;
  wire \nand_12.nand_2 ;
  wire \nand_12.nand_3 ;
  wire \nand_12.nand_4 ;
  wire \nand_12.out ;
  wire \nand_13.and_0 ;
  wire \nand_13.and_1 ;
  wire \nand_13.and_2 ;
  wire \nand_13.and_3 ;
  wire \nand_13.and_4 ;
  wire \nand_13.in_0 ;
  wire \nand_13.in_1 ;
  wire \nand_13.in_2 ;
  wire \nand_13.in_3 ;
  wire \nand_13.in_4 ;
  wire \nand_13.in_5 ;
  wire \nand_13.in_6 ;
  wire \nand_13.nand_0 ;
  wire \nand_13.nand_1 ;
  wire \nand_13.nand_2 ;
  wire \nand_13.nand_3 ;
  wire \nand_13.nand_4 ;
  wire \nand_13.out ;
  wire \nand_14.and_0 ;
  wire \nand_14.and_1 ;
  wire \nand_14.and_2 ;
  wire \nand_14.and_3 ;
  wire \nand_14.and_4 ;
  wire \nand_14.in_0 ;
  wire \nand_14.in_1 ;
  wire \nand_14.in_2 ;
  wire \nand_14.in_3 ;
  wire \nand_14.in_4 ;
  wire \nand_14.in_5 ;
  wire \nand_14.in_6 ;
  wire \nand_14.nand_0 ;
  wire \nand_14.nand_1 ;
  wire \nand_14.nand_2 ;
  wire \nand_14.nand_3 ;
  wire \nand_14.nand_4 ;
  wire \nand_14.out ;
  wire \nand_15.and_0 ;
  wire \nand_15.and_1 ;
  wire \nand_15.and_2 ;
  wire \nand_15.and_3 ;
  wire \nand_15.and_4 ;
  wire \nand_15.in_0 ;
  wire \nand_15.in_1 ;
  wire \nand_15.in_2 ;
  wire \nand_15.in_3 ;
  wire \nand_15.in_4 ;
  wire \nand_15.in_5 ;
  wire \nand_15.in_6 ;
  wire \nand_15.nand_0 ;
  wire \nand_15.nand_1 ;
  wire \nand_15.nand_2 ;
  wire \nand_15.nand_3 ;
  wire \nand_15.nand_4 ;
  wire \nand_15.out ;
  wire \nand_16.and_0 ;
  wire \nand_16.and_1 ;
  wire \nand_16.and_2 ;
  wire \nand_16.and_3 ;
  wire \nand_16.and_4 ;
  wire \nand_16.in_0 ;
  wire \nand_16.in_1 ;
  wire \nand_16.in_2 ;
  wire \nand_16.in_3 ;
  wire \nand_16.in_4 ;
  wire \nand_16.in_5 ;
  wire \nand_16.in_6 ;
  wire \nand_16.nand_0 ;
  wire \nand_16.nand_1 ;
  wire \nand_16.nand_2 ;
  wire \nand_16.nand_3 ;
  wire \nand_16.nand_4 ;
  wire \nand_16.out ;
  wire \nand_17.and_0 ;
  wire \nand_17.and_1 ;
  wire \nand_17.and_2 ;
  wire \nand_17.and_3 ;
  wire \nand_17.and_4 ;
  wire \nand_17.in_0 ;
  wire \nand_17.in_1 ;
  wire \nand_17.in_2 ;
  wire \nand_17.in_3 ;
  wire \nand_17.in_4 ;
  wire \nand_17.in_5 ;
  wire \nand_17.in_6 ;
  wire \nand_17.nand_0 ;
  wire \nand_17.nand_1 ;
  wire \nand_17.nand_2 ;
  wire \nand_17.nand_3 ;
  wire \nand_17.nand_4 ;
  wire \nand_17.out ;
  wire \nand_18.and_0 ;
  wire \nand_18.and_1 ;
  wire \nand_18.and_2 ;
  wire \nand_18.and_3 ;
  wire \nand_18.and_4 ;
  wire \nand_18.in_0 ;
  wire \nand_18.in_1 ;
  wire \nand_18.in_2 ;
  wire \nand_18.in_3 ;
  wire \nand_18.in_4 ;
  wire \nand_18.in_5 ;
  wire \nand_18.in_6 ;
  wire \nand_18.nand_0 ;
  wire \nand_18.nand_1 ;
  wire \nand_18.nand_2 ;
  wire \nand_18.nand_3 ;
  wire \nand_18.nand_4 ;
  wire \nand_18.out ;
  wire \nand_19.and_0 ;
  wire \nand_19.and_1 ;
  wire \nand_19.and_2 ;
  wire \nand_19.and_3 ;
  wire \nand_19.and_4 ;
  wire \nand_19.in_0 ;
  wire \nand_19.in_1 ;
  wire \nand_19.in_2 ;
  wire \nand_19.in_3 ;
  wire \nand_19.in_4 ;
  wire \nand_19.in_5 ;
  wire \nand_19.in_6 ;
  wire \nand_19.nand_0 ;
  wire \nand_19.nand_1 ;
  wire \nand_19.nand_2 ;
  wire \nand_19.nand_3 ;
  wire \nand_19.nand_4 ;
  wire \nand_19.out ;
  wire \nand_2.and_0 ;
  wire \nand_2.and_1 ;
  wire \nand_2.and_2 ;
  wire \nand_2.and_3 ;
  wire \nand_2.and_4 ;
  wire \nand_2.in_0 ;
  wire \nand_2.in_1 ;
  wire \nand_2.in_2 ;
  wire \nand_2.in_3 ;
  wire \nand_2.in_4 ;
  wire \nand_2.in_5 ;
  wire \nand_2.in_6 ;
  wire \nand_2.nand_0 ;
  wire \nand_2.nand_1 ;
  wire \nand_2.nand_2 ;
  wire \nand_2.nand_3 ;
  wire \nand_2.nand_4 ;
  wire \nand_2.out ;
  wire \nand_20.and_0 ;
  wire \nand_20.and_1 ;
  wire \nand_20.and_2 ;
  wire \nand_20.and_3 ;
  wire \nand_20.and_4 ;
  wire \nand_20.in_0 ;
  wire \nand_20.in_1 ;
  wire \nand_20.in_2 ;
  wire \nand_20.in_3 ;
  wire \nand_20.in_4 ;
  wire \nand_20.in_5 ;
  wire \nand_20.in_6 ;
  wire \nand_20.nand_0 ;
  wire \nand_20.nand_1 ;
  wire \nand_20.nand_2 ;
  wire \nand_20.nand_3 ;
  wire \nand_20.nand_4 ;
  wire \nand_20.out ;
  wire \nand_21.and_0 ;
  wire \nand_21.and_1 ;
  wire \nand_21.and_2 ;
  wire \nand_21.and_3 ;
  wire \nand_21.and_4 ;
  wire \nand_21.in_0 ;
  wire \nand_21.in_1 ;
  wire \nand_21.in_2 ;
  wire \nand_21.in_3 ;
  wire \nand_21.in_4 ;
  wire \nand_21.in_5 ;
  wire \nand_21.in_6 ;
  wire \nand_21.nand_0 ;
  wire \nand_21.nand_1 ;
  wire \nand_21.nand_2 ;
  wire \nand_21.nand_3 ;
  wire \nand_21.nand_4 ;
  wire \nand_21.out ;
  wire \nand_22.and_0 ;
  wire \nand_22.and_1 ;
  wire \nand_22.and_2 ;
  wire \nand_22.and_3 ;
  wire \nand_22.and_4 ;
  wire \nand_22.in_0 ;
  wire \nand_22.in_1 ;
  wire \nand_22.in_2 ;
  wire \nand_22.in_3 ;
  wire \nand_22.in_4 ;
  wire \nand_22.in_5 ;
  wire \nand_22.in_6 ;
  wire \nand_22.nand_0 ;
  wire \nand_22.nand_1 ;
  wire \nand_22.nand_2 ;
  wire \nand_22.nand_3 ;
  wire \nand_22.nand_4 ;
  wire \nand_22.out ;
  wire \nand_23.and_0 ;
  wire \nand_23.and_1 ;
  wire \nand_23.and_2 ;
  wire \nand_23.and_3 ;
  wire \nand_23.and_4 ;
  wire \nand_23.in_0 ;
  wire \nand_23.in_1 ;
  wire \nand_23.in_2 ;
  wire \nand_23.in_3 ;
  wire \nand_23.in_4 ;
  wire \nand_23.in_5 ;
  wire \nand_23.in_6 ;
  wire \nand_23.nand_0 ;
  wire \nand_23.nand_1 ;
  wire \nand_23.nand_2 ;
  wire \nand_23.nand_3 ;
  wire \nand_23.nand_4 ;
  wire \nand_23.out ;
  wire \nand_24.and_0 ;
  wire \nand_24.and_1 ;
  wire \nand_24.and_2 ;
  wire \nand_24.and_3 ;
  wire \nand_24.and_4 ;
  wire \nand_24.in_0 ;
  wire \nand_24.in_1 ;
  wire \nand_24.in_2 ;
  wire \nand_24.in_3 ;
  wire \nand_24.in_4 ;
  wire \nand_24.in_5 ;
  wire \nand_24.in_6 ;
  wire \nand_24.nand_0 ;
  wire \nand_24.nand_1 ;
  wire \nand_24.nand_2 ;
  wire \nand_24.nand_3 ;
  wire \nand_24.nand_4 ;
  wire \nand_24.out ;
  wire \nand_25.and_0 ;
  wire \nand_25.and_1 ;
  wire \nand_25.and_2 ;
  wire \nand_25.and_3 ;
  wire \nand_25.and_4 ;
  wire \nand_25.in_0 ;
  wire \nand_25.in_1 ;
  wire \nand_25.in_2 ;
  wire \nand_25.in_3 ;
  wire \nand_25.in_4 ;
  wire \nand_25.in_5 ;
  wire \nand_25.in_6 ;
  wire \nand_25.nand_0 ;
  wire \nand_25.nand_1 ;
  wire \nand_25.nand_2 ;
  wire \nand_25.nand_3 ;
  wire \nand_25.nand_4 ;
  wire \nand_25.out ;
  wire \nand_26.and_0 ;
  wire \nand_26.and_1 ;
  wire \nand_26.and_2 ;
  wire \nand_26.and_3 ;
  wire \nand_26.and_4 ;
  wire \nand_26.in_0 ;
  wire \nand_26.in_1 ;
  wire \nand_26.in_2 ;
  wire \nand_26.in_3 ;
  wire \nand_26.in_4 ;
  wire \nand_26.in_5 ;
  wire \nand_26.in_6 ;
  wire \nand_26.nand_0 ;
  wire \nand_26.nand_1 ;
  wire \nand_26.nand_2 ;
  wire \nand_26.nand_3 ;
  wire \nand_26.nand_4 ;
  wire \nand_26.out ;
  wire \nand_27.and_0 ;
  wire \nand_27.and_1 ;
  wire \nand_27.and_2 ;
  wire \nand_27.and_3 ;
  wire \nand_27.and_4 ;
  wire \nand_27.in_0 ;
  wire \nand_27.in_1 ;
  wire \nand_27.in_2 ;
  wire \nand_27.in_3 ;
  wire \nand_27.in_4 ;
  wire \nand_27.in_5 ;
  wire \nand_27.in_6 ;
  wire \nand_27.nand_0 ;
  wire \nand_27.nand_1 ;
  wire \nand_27.nand_2 ;
  wire \nand_27.nand_3 ;
  wire \nand_27.nand_4 ;
  wire \nand_27.out ;
  wire \nand_28.and_0 ;
  wire \nand_28.and_1 ;
  wire \nand_28.and_2 ;
  wire \nand_28.and_3 ;
  wire \nand_28.and_4 ;
  wire \nand_28.in_0 ;
  wire \nand_28.in_1 ;
  wire \nand_28.in_2 ;
  wire \nand_28.in_3 ;
  wire \nand_28.in_4 ;
  wire \nand_28.in_5 ;
  wire \nand_28.in_6 ;
  wire \nand_28.nand_0 ;
  wire \nand_28.nand_1 ;
  wire \nand_28.nand_2 ;
  wire \nand_28.nand_3 ;
  wire \nand_28.nand_4 ;
  wire \nand_28.out ;
  wire \nand_29.and_0 ;
  wire \nand_29.and_1 ;
  wire \nand_29.and_2 ;
  wire \nand_29.and_3 ;
  wire \nand_29.and_4 ;
  wire \nand_29.in_0 ;
  wire \nand_29.in_1 ;
  wire \nand_29.in_2 ;
  wire \nand_29.in_3 ;
  wire \nand_29.in_4 ;
  wire \nand_29.in_5 ;
  wire \nand_29.in_6 ;
  wire \nand_29.nand_0 ;
  wire \nand_29.nand_1 ;
  wire \nand_29.nand_2 ;
  wire \nand_29.nand_3 ;
  wire \nand_29.nand_4 ;
  wire \nand_29.out ;
  wire \nand_3.and_0 ;
  wire \nand_3.and_1 ;
  wire \nand_3.and_2 ;
  wire \nand_3.and_3 ;
  wire \nand_3.and_4 ;
  wire \nand_3.in_0 ;
  wire \nand_3.in_1 ;
  wire \nand_3.in_2 ;
  wire \nand_3.in_3 ;
  wire \nand_3.in_4 ;
  wire \nand_3.in_5 ;
  wire \nand_3.in_6 ;
  wire \nand_3.nand_0 ;
  wire \nand_3.nand_1 ;
  wire \nand_3.nand_2 ;
  wire \nand_3.nand_3 ;
  wire \nand_3.nand_4 ;
  wire \nand_3.out ;
  wire \nand_30.and_0 ;
  wire \nand_30.and_1 ;
  wire \nand_30.and_2 ;
  wire \nand_30.and_3 ;
  wire \nand_30.and_4 ;
  wire \nand_30.in_0 ;
  wire \nand_30.in_1 ;
  wire \nand_30.in_2 ;
  wire \nand_30.in_3 ;
  wire \nand_30.in_4 ;
  wire \nand_30.in_5 ;
  wire \nand_30.in_6 ;
  wire \nand_30.nand_0 ;
  wire \nand_30.nand_1 ;
  wire \nand_30.nand_2 ;
  wire \nand_30.nand_3 ;
  wire \nand_30.nand_4 ;
  wire \nand_30.out ;
  wire \nand_31.and_0 ;
  wire \nand_31.and_1 ;
  wire \nand_31.and_2 ;
  wire \nand_31.and_3 ;
  wire \nand_31.and_4 ;
  wire \nand_31.in_0 ;
  wire \nand_31.in_1 ;
  wire \nand_31.in_2 ;
  wire \nand_31.in_3 ;
  wire \nand_31.in_4 ;
  wire \nand_31.in_5 ;
  wire \nand_31.in_6 ;
  wire \nand_31.nand_0 ;
  wire \nand_31.nand_1 ;
  wire \nand_31.nand_2 ;
  wire \nand_31.nand_3 ;
  wire \nand_31.nand_4 ;
  wire \nand_31.out ;
  wire \nand_32.and_0 ;
  wire \nand_32.and_1 ;
  wire \nand_32.and_2 ;
  wire \nand_32.and_3 ;
  wire \nand_32.and_4 ;
  wire \nand_32.in_0 ;
  wire \nand_32.in_1 ;
  wire \nand_32.in_2 ;
  wire \nand_32.in_3 ;
  wire \nand_32.in_4 ;
  wire \nand_32.in_5 ;
  wire \nand_32.in_6 ;
  wire \nand_32.nand_0 ;
  wire \nand_32.nand_1 ;
  wire \nand_32.nand_2 ;
  wire \nand_32.nand_3 ;
  wire \nand_32.nand_4 ;
  wire \nand_32.out ;
  wire \nand_33.and_0 ;
  wire \nand_33.and_1 ;
  wire \nand_33.and_2 ;
  wire \nand_33.and_3 ;
  wire \nand_33.and_4 ;
  wire \nand_33.in_0 ;
  wire \nand_33.in_1 ;
  wire \nand_33.in_2 ;
  wire \nand_33.in_3 ;
  wire \nand_33.in_4 ;
  wire \nand_33.in_5 ;
  wire \nand_33.in_6 ;
  wire \nand_33.nand_0 ;
  wire \nand_33.nand_1 ;
  wire \nand_33.nand_2 ;
  wire \nand_33.nand_3 ;
  wire \nand_33.nand_4 ;
  wire \nand_33.out ;
  wire \nand_34.and_0 ;
  wire \nand_34.and_1 ;
  wire \nand_34.and_2 ;
  wire \nand_34.and_3 ;
  wire \nand_34.and_4 ;
  wire \nand_34.in_0 ;
  wire \nand_34.in_1 ;
  wire \nand_34.in_2 ;
  wire \nand_34.in_3 ;
  wire \nand_34.in_4 ;
  wire \nand_34.in_5 ;
  wire \nand_34.in_6 ;
  wire \nand_34.nand_0 ;
  wire \nand_34.nand_1 ;
  wire \nand_34.nand_2 ;
  wire \nand_34.nand_3 ;
  wire \nand_34.nand_4 ;
  wire \nand_34.out ;
  wire \nand_35.and_0 ;
  wire \nand_35.and_1 ;
  wire \nand_35.and_2 ;
  wire \nand_35.and_3 ;
  wire \nand_35.and_4 ;
  wire \nand_35.in_0 ;
  wire \nand_35.in_1 ;
  wire \nand_35.in_2 ;
  wire \nand_35.in_3 ;
  wire \nand_35.in_4 ;
  wire \nand_35.in_5 ;
  wire \nand_35.in_6 ;
  wire \nand_35.nand_0 ;
  wire \nand_35.nand_1 ;
  wire \nand_35.nand_2 ;
  wire \nand_35.nand_3 ;
  wire \nand_35.nand_4 ;
  wire \nand_35.out ;
  wire \nand_36.and_0 ;
  wire \nand_36.and_1 ;
  wire \nand_36.and_2 ;
  wire \nand_36.and_3 ;
  wire \nand_36.and_4 ;
  wire \nand_36.in_0 ;
  wire \nand_36.in_1 ;
  wire \nand_36.in_2 ;
  wire \nand_36.in_3 ;
  wire \nand_36.in_4 ;
  wire \nand_36.in_5 ;
  wire \nand_36.in_6 ;
  wire \nand_36.nand_0 ;
  wire \nand_36.nand_1 ;
  wire \nand_36.nand_2 ;
  wire \nand_36.nand_3 ;
  wire \nand_36.nand_4 ;
  wire \nand_36.out ;
  wire \nand_37.and_0 ;
  wire \nand_37.and_1 ;
  wire \nand_37.and_2 ;
  wire \nand_37.and_3 ;
  wire \nand_37.and_4 ;
  wire \nand_37.in_0 ;
  wire \nand_37.in_1 ;
  wire \nand_37.in_2 ;
  wire \nand_37.in_3 ;
  wire \nand_37.in_4 ;
  wire \nand_37.in_5 ;
  wire \nand_37.in_6 ;
  wire \nand_37.nand_0 ;
  wire \nand_37.nand_1 ;
  wire \nand_37.nand_2 ;
  wire \nand_37.nand_3 ;
  wire \nand_37.nand_4 ;
  wire \nand_37.out ;
  wire \nand_38.and_0 ;
  wire \nand_38.and_1 ;
  wire \nand_38.and_2 ;
  wire \nand_38.and_3 ;
  wire \nand_38.and_4 ;
  wire \nand_38.in_0 ;
  wire \nand_38.in_1 ;
  wire \nand_38.in_2 ;
  wire \nand_38.in_3 ;
  wire \nand_38.in_4 ;
  wire \nand_38.in_5 ;
  wire \nand_38.in_6 ;
  wire \nand_38.nand_0 ;
  wire \nand_38.nand_1 ;
  wire \nand_38.nand_2 ;
  wire \nand_38.nand_3 ;
  wire \nand_38.nand_4 ;
  wire \nand_38.out ;
  wire \nand_39.and_0 ;
  wire \nand_39.and_1 ;
  wire \nand_39.and_2 ;
  wire \nand_39.and_3 ;
  wire \nand_39.and_4 ;
  wire \nand_39.in_0 ;
  wire \nand_39.in_1 ;
  wire \nand_39.in_2 ;
  wire \nand_39.in_3 ;
  wire \nand_39.in_4 ;
  wire \nand_39.in_5 ;
  wire \nand_39.in_6 ;
  wire \nand_39.nand_0 ;
  wire \nand_39.nand_1 ;
  wire \nand_39.nand_2 ;
  wire \nand_39.nand_3 ;
  wire \nand_39.nand_4 ;
  wire \nand_39.out ;
  wire \nand_4.and_0 ;
  wire \nand_4.and_1 ;
  wire \nand_4.and_2 ;
  wire \nand_4.and_3 ;
  wire \nand_4.and_4 ;
  wire \nand_4.in_0 ;
  wire \nand_4.in_1 ;
  wire \nand_4.in_2 ;
  wire \nand_4.in_3 ;
  wire \nand_4.in_4 ;
  wire \nand_4.in_5 ;
  wire \nand_4.in_6 ;
  wire \nand_4.nand_0 ;
  wire \nand_4.nand_1 ;
  wire \nand_4.nand_2 ;
  wire \nand_4.nand_3 ;
  wire \nand_4.nand_4 ;
  wire \nand_4.out ;
  wire \nand_40.and_0 ;
  wire \nand_40.and_1 ;
  wire \nand_40.and_2 ;
  wire \nand_40.and_3 ;
  wire \nand_40.and_4 ;
  wire \nand_40.in_0 ;
  wire \nand_40.in_1 ;
  wire \nand_40.in_2 ;
  wire \nand_40.in_3 ;
  wire \nand_40.in_4 ;
  wire \nand_40.in_5 ;
  wire \nand_40.in_6 ;
  wire \nand_40.nand_0 ;
  wire \nand_40.nand_1 ;
  wire \nand_40.nand_2 ;
  wire \nand_40.nand_3 ;
  wire \nand_40.nand_4 ;
  wire \nand_40.out ;
  wire \nand_41.and_0 ;
  wire \nand_41.and_1 ;
  wire \nand_41.and_2 ;
  wire \nand_41.and_3 ;
  wire \nand_41.and_4 ;
  wire \nand_41.in_0 ;
  wire \nand_41.in_1 ;
  wire \nand_41.in_2 ;
  wire \nand_41.in_3 ;
  wire \nand_41.in_4 ;
  wire \nand_41.in_5 ;
  wire \nand_41.in_6 ;
  wire \nand_41.nand_0 ;
  wire \nand_41.nand_1 ;
  wire \nand_41.nand_2 ;
  wire \nand_41.nand_3 ;
  wire \nand_41.nand_4 ;
  wire \nand_41.out ;
  wire \nand_42.and_0 ;
  wire \nand_42.and_1 ;
  wire \nand_42.and_2 ;
  wire \nand_42.and_3 ;
  wire \nand_42.and_4 ;
  wire \nand_42.in_0 ;
  wire \nand_42.in_1 ;
  wire \nand_42.in_2 ;
  wire \nand_42.in_3 ;
  wire \nand_42.in_4 ;
  wire \nand_42.in_5 ;
  wire \nand_42.in_6 ;
  wire \nand_42.nand_0 ;
  wire \nand_42.nand_1 ;
  wire \nand_42.nand_2 ;
  wire \nand_42.nand_3 ;
  wire \nand_42.nand_4 ;
  wire \nand_42.out ;
  wire \nand_43.and_0 ;
  wire \nand_43.and_1 ;
  wire \nand_43.and_2 ;
  wire \nand_43.and_3 ;
  wire \nand_43.and_4 ;
  wire \nand_43.in_0 ;
  wire \nand_43.in_1 ;
  wire \nand_43.in_2 ;
  wire \nand_43.in_3 ;
  wire \nand_43.in_4 ;
  wire \nand_43.in_5 ;
  wire \nand_43.in_6 ;
  wire \nand_43.nand_0 ;
  wire \nand_43.nand_1 ;
  wire \nand_43.nand_2 ;
  wire \nand_43.nand_3 ;
  wire \nand_43.nand_4 ;
  wire \nand_43.out ;
  wire \nand_44.and_0 ;
  wire \nand_44.and_1 ;
  wire \nand_44.and_2 ;
  wire \nand_44.and_3 ;
  wire \nand_44.and_4 ;
  wire \nand_44.in_0 ;
  wire \nand_44.in_1 ;
  wire \nand_44.in_2 ;
  wire \nand_44.in_3 ;
  wire \nand_44.in_4 ;
  wire \nand_44.in_5 ;
  wire \nand_44.in_6 ;
  wire \nand_44.nand_0 ;
  wire \nand_44.nand_1 ;
  wire \nand_44.nand_2 ;
  wire \nand_44.nand_3 ;
  wire \nand_44.nand_4 ;
  wire \nand_44.out ;
  wire \nand_45.and_0 ;
  wire \nand_45.and_1 ;
  wire \nand_45.and_2 ;
  wire \nand_45.and_3 ;
  wire \nand_45.and_4 ;
  wire \nand_45.in_0 ;
  wire \nand_45.in_1 ;
  wire \nand_45.in_2 ;
  wire \nand_45.in_3 ;
  wire \nand_45.in_4 ;
  wire \nand_45.in_5 ;
  wire \nand_45.in_6 ;
  wire \nand_45.nand_0 ;
  wire \nand_45.nand_1 ;
  wire \nand_45.nand_2 ;
  wire \nand_45.nand_3 ;
  wire \nand_45.nand_4 ;
  wire \nand_45.out ;
  wire \nand_46.and_0 ;
  wire \nand_46.and_1 ;
  wire \nand_46.and_2 ;
  wire \nand_46.and_3 ;
  wire \nand_46.and_4 ;
  wire \nand_46.in_0 ;
  wire \nand_46.in_1 ;
  wire \nand_46.in_2 ;
  wire \nand_46.in_3 ;
  wire \nand_46.in_4 ;
  wire \nand_46.in_5 ;
  wire \nand_46.in_6 ;
  wire \nand_46.nand_0 ;
  wire \nand_46.nand_1 ;
  wire \nand_46.nand_2 ;
  wire \nand_46.nand_3 ;
  wire \nand_46.nand_4 ;
  wire \nand_46.out ;
  wire \nand_47.and_0 ;
  wire \nand_47.and_1 ;
  wire \nand_47.and_2 ;
  wire \nand_47.and_3 ;
  wire \nand_47.and_4 ;
  wire \nand_47.in_0 ;
  wire \nand_47.in_1 ;
  wire \nand_47.in_2 ;
  wire \nand_47.in_3 ;
  wire \nand_47.in_4 ;
  wire \nand_47.in_5 ;
  wire \nand_47.in_6 ;
  wire \nand_47.nand_0 ;
  wire \nand_47.nand_1 ;
  wire \nand_47.nand_2 ;
  wire \nand_47.nand_3 ;
  wire \nand_47.nand_4 ;
  wire \nand_47.out ;
  wire \nand_48.and_0 ;
  wire \nand_48.and_1 ;
  wire \nand_48.and_2 ;
  wire \nand_48.and_3 ;
  wire \nand_48.and_4 ;
  wire \nand_48.in_0 ;
  wire \nand_48.in_1 ;
  wire \nand_48.in_2 ;
  wire \nand_48.in_3 ;
  wire \nand_48.in_4 ;
  wire \nand_48.in_5 ;
  wire \nand_48.in_6 ;
  wire \nand_48.nand_0 ;
  wire \nand_48.nand_1 ;
  wire \nand_48.nand_2 ;
  wire \nand_48.nand_3 ;
  wire \nand_48.nand_4 ;
  wire \nand_48.out ;
  wire \nand_49.and_0 ;
  wire \nand_49.and_1 ;
  wire \nand_49.and_2 ;
  wire \nand_49.and_3 ;
  wire \nand_49.and_4 ;
  wire \nand_49.in_0 ;
  wire \nand_49.in_1 ;
  wire \nand_49.in_2 ;
  wire \nand_49.in_3 ;
  wire \nand_49.in_4 ;
  wire \nand_49.in_5 ;
  wire \nand_49.in_6 ;
  wire \nand_49.nand_0 ;
  wire \nand_49.nand_1 ;
  wire \nand_49.nand_2 ;
  wire \nand_49.nand_3 ;
  wire \nand_49.nand_4 ;
  wire \nand_49.out ;
  wire \nand_5.and_0 ;
  wire \nand_5.and_1 ;
  wire \nand_5.and_2 ;
  wire \nand_5.and_3 ;
  wire \nand_5.and_4 ;
  wire \nand_5.in_0 ;
  wire \nand_5.in_1 ;
  wire \nand_5.in_2 ;
  wire \nand_5.in_3 ;
  wire \nand_5.in_4 ;
  wire \nand_5.in_5 ;
  wire \nand_5.in_6 ;
  wire \nand_5.nand_0 ;
  wire \nand_5.nand_1 ;
  wire \nand_5.nand_2 ;
  wire \nand_5.nand_3 ;
  wire \nand_5.nand_4 ;
  wire \nand_5.out ;
  wire \nand_50.and_0 ;
  wire \nand_50.and_1 ;
  wire \nand_50.and_2 ;
  wire \nand_50.and_3 ;
  wire \nand_50.and_4 ;
  wire \nand_50.in_0 ;
  wire \nand_50.in_1 ;
  wire \nand_50.in_2 ;
  wire \nand_50.in_3 ;
  wire \nand_50.in_4 ;
  wire \nand_50.in_5 ;
  wire \nand_50.in_6 ;
  wire \nand_50.nand_0 ;
  wire \nand_50.nand_1 ;
  wire \nand_50.nand_2 ;
  wire \nand_50.nand_3 ;
  wire \nand_50.nand_4 ;
  wire \nand_50.out ;
  wire \nand_51.and_0 ;
  wire \nand_51.and_1 ;
  wire \nand_51.and_2 ;
  wire \nand_51.and_3 ;
  wire \nand_51.and_4 ;
  wire \nand_51.in_0 ;
  wire \nand_51.in_1 ;
  wire \nand_51.in_2 ;
  wire \nand_51.in_3 ;
  wire \nand_51.in_4 ;
  wire \nand_51.in_5 ;
  wire \nand_51.in_6 ;
  wire \nand_51.nand_0 ;
  wire \nand_51.nand_1 ;
  wire \nand_51.nand_2 ;
  wire \nand_51.nand_3 ;
  wire \nand_51.nand_4 ;
  wire \nand_51.out ;
  wire \nand_52.and_0 ;
  wire \nand_52.and_1 ;
  wire \nand_52.and_2 ;
  wire \nand_52.and_3 ;
  wire \nand_52.and_4 ;
  wire \nand_52.in_0 ;
  wire \nand_52.in_1 ;
  wire \nand_52.in_2 ;
  wire \nand_52.in_3 ;
  wire \nand_52.in_4 ;
  wire \nand_52.in_5 ;
  wire \nand_52.in_6 ;
  wire \nand_52.nand_0 ;
  wire \nand_52.nand_1 ;
  wire \nand_52.nand_2 ;
  wire \nand_52.nand_3 ;
  wire \nand_52.nand_4 ;
  wire \nand_52.out ;
  wire \nand_53.and_0 ;
  wire \nand_53.and_1 ;
  wire \nand_53.and_2 ;
  wire \nand_53.and_3 ;
  wire \nand_53.and_4 ;
  wire \nand_53.in_0 ;
  wire \nand_53.in_1 ;
  wire \nand_53.in_2 ;
  wire \nand_53.in_3 ;
  wire \nand_53.in_4 ;
  wire \nand_53.in_5 ;
  wire \nand_53.in_6 ;
  wire \nand_53.nand_0 ;
  wire \nand_53.nand_1 ;
  wire \nand_53.nand_2 ;
  wire \nand_53.nand_3 ;
  wire \nand_53.nand_4 ;
  wire \nand_53.out ;
  wire \nand_54.and_0 ;
  wire \nand_54.and_1 ;
  wire \nand_54.and_2 ;
  wire \nand_54.and_3 ;
  wire \nand_54.and_4 ;
  wire \nand_54.in_0 ;
  wire \nand_54.in_1 ;
  wire \nand_54.in_2 ;
  wire \nand_54.in_3 ;
  wire \nand_54.in_4 ;
  wire \nand_54.in_5 ;
  wire \nand_54.in_6 ;
  wire \nand_54.nand_0 ;
  wire \nand_54.nand_1 ;
  wire \nand_54.nand_2 ;
  wire \nand_54.nand_3 ;
  wire \nand_54.nand_4 ;
  wire \nand_54.out ;
  wire \nand_55.and_0 ;
  wire \nand_55.and_1 ;
  wire \nand_55.and_2 ;
  wire \nand_55.and_3 ;
  wire \nand_55.and_4 ;
  wire \nand_55.in_0 ;
  wire \nand_55.in_1 ;
  wire \nand_55.in_2 ;
  wire \nand_55.in_3 ;
  wire \nand_55.in_4 ;
  wire \nand_55.in_5 ;
  wire \nand_55.in_6 ;
  wire \nand_55.nand_0 ;
  wire \nand_55.nand_1 ;
  wire \nand_55.nand_2 ;
  wire \nand_55.nand_3 ;
  wire \nand_55.nand_4 ;
  wire \nand_55.out ;
  wire \nand_56.and_0 ;
  wire \nand_56.and_1 ;
  wire \nand_56.and_2 ;
  wire \nand_56.and_3 ;
  wire \nand_56.and_4 ;
  wire \nand_56.in_0 ;
  wire \nand_56.in_1 ;
  wire \nand_56.in_2 ;
  wire \nand_56.in_3 ;
  wire \nand_56.in_4 ;
  wire \nand_56.in_5 ;
  wire \nand_56.in_6 ;
  wire \nand_56.nand_0 ;
  wire \nand_56.nand_1 ;
  wire \nand_56.nand_2 ;
  wire \nand_56.nand_3 ;
  wire \nand_56.nand_4 ;
  wire \nand_56.out ;
  wire \nand_57.and_0 ;
  wire \nand_57.and_1 ;
  wire \nand_57.and_2 ;
  wire \nand_57.and_3 ;
  wire \nand_57.and_4 ;
  wire \nand_57.in_0 ;
  wire \nand_57.in_1 ;
  wire \nand_57.in_2 ;
  wire \nand_57.in_3 ;
  wire \nand_57.in_4 ;
  wire \nand_57.in_5 ;
  wire \nand_57.in_6 ;
  wire \nand_57.nand_0 ;
  wire \nand_57.nand_1 ;
  wire \nand_57.nand_2 ;
  wire \nand_57.nand_3 ;
  wire \nand_57.nand_4 ;
  wire \nand_57.out ;
  wire \nand_58.and_0 ;
  wire \nand_58.and_1 ;
  wire \nand_58.and_2 ;
  wire \nand_58.and_3 ;
  wire \nand_58.and_4 ;
  wire \nand_58.in_0 ;
  wire \nand_58.in_1 ;
  wire \nand_58.in_2 ;
  wire \nand_58.in_3 ;
  wire \nand_58.in_4 ;
  wire \nand_58.in_5 ;
  wire \nand_58.in_6 ;
  wire \nand_58.nand_0 ;
  wire \nand_58.nand_1 ;
  wire \nand_58.nand_2 ;
  wire \nand_58.nand_3 ;
  wire \nand_58.nand_4 ;
  wire \nand_58.out ;
  wire \nand_59.and_0 ;
  wire \nand_59.and_1 ;
  wire \nand_59.and_2 ;
  wire \nand_59.and_3 ;
  wire \nand_59.and_4 ;
  wire \nand_59.in_0 ;
  wire \nand_59.in_1 ;
  wire \nand_59.in_2 ;
  wire \nand_59.in_3 ;
  wire \nand_59.in_4 ;
  wire \nand_59.in_5 ;
  wire \nand_59.in_6 ;
  wire \nand_59.nand_0 ;
  wire \nand_59.nand_1 ;
  wire \nand_59.nand_2 ;
  wire \nand_59.nand_3 ;
  wire \nand_59.nand_4 ;
  wire \nand_59.out ;
  wire \nand_6.and_0 ;
  wire \nand_6.and_1 ;
  wire \nand_6.and_2 ;
  wire \nand_6.and_3 ;
  wire \nand_6.and_4 ;
  wire \nand_6.in_0 ;
  wire \nand_6.in_1 ;
  wire \nand_6.in_2 ;
  wire \nand_6.in_3 ;
  wire \nand_6.in_4 ;
  wire \nand_6.in_5 ;
  wire \nand_6.in_6 ;
  wire \nand_6.nand_0 ;
  wire \nand_6.nand_1 ;
  wire \nand_6.nand_2 ;
  wire \nand_6.nand_3 ;
  wire \nand_6.nand_4 ;
  wire \nand_6.out ;
  wire \nand_60.and_0 ;
  wire \nand_60.and_1 ;
  wire \nand_60.and_2 ;
  wire \nand_60.and_3 ;
  wire \nand_60.and_4 ;
  wire \nand_60.in_0 ;
  wire \nand_60.in_1 ;
  wire \nand_60.in_2 ;
  wire \nand_60.in_3 ;
  wire \nand_60.in_4 ;
  wire \nand_60.in_5 ;
  wire \nand_60.in_6 ;
  wire \nand_60.nand_0 ;
  wire \nand_60.nand_1 ;
  wire \nand_60.nand_2 ;
  wire \nand_60.nand_3 ;
  wire \nand_60.nand_4 ;
  wire \nand_60.out ;
  wire \nand_61.and_0 ;
  wire \nand_61.and_1 ;
  wire \nand_61.and_2 ;
  wire \nand_61.and_3 ;
  wire \nand_61.and_4 ;
  wire \nand_61.in_0 ;
  wire \nand_61.in_1 ;
  wire \nand_61.in_2 ;
  wire \nand_61.in_3 ;
  wire \nand_61.in_4 ;
  wire \nand_61.in_5 ;
  wire \nand_61.in_6 ;
  wire \nand_61.nand_0 ;
  wire \nand_61.nand_1 ;
  wire \nand_61.nand_2 ;
  wire \nand_61.nand_3 ;
  wire \nand_61.nand_4 ;
  wire \nand_61.out ;
  wire \nand_62.and_0 ;
  wire \nand_62.and_1 ;
  wire \nand_62.and_2 ;
  wire \nand_62.and_3 ;
  wire \nand_62.and_4 ;
  wire \nand_62.in_0 ;
  wire \nand_62.in_1 ;
  wire \nand_62.in_2 ;
  wire \nand_62.in_3 ;
  wire \nand_62.in_4 ;
  wire \nand_62.in_5 ;
  wire \nand_62.in_6 ;
  wire \nand_62.nand_0 ;
  wire \nand_62.nand_1 ;
  wire \nand_62.nand_2 ;
  wire \nand_62.nand_3 ;
  wire \nand_62.nand_4 ;
  wire \nand_62.out ;
  wire \nand_63.and_0 ;
  wire \nand_63.and_1 ;
  wire \nand_63.and_2 ;
  wire \nand_63.and_3 ;
  wire \nand_63.and_4 ;
  wire \nand_63.in_0 ;
  wire \nand_63.in_1 ;
  wire \nand_63.in_2 ;
  wire \nand_63.in_3 ;
  wire \nand_63.in_4 ;
  wire \nand_63.in_5 ;
  wire \nand_63.in_6 ;
  wire \nand_63.nand_0 ;
  wire \nand_63.nand_1 ;
  wire \nand_63.nand_2 ;
  wire \nand_63.nand_3 ;
  wire \nand_63.nand_4 ;
  wire \nand_63.out ;
  wire \nand_7.and_0 ;
  wire \nand_7.and_1 ;
  wire \nand_7.and_2 ;
  wire \nand_7.and_3 ;
  wire \nand_7.and_4 ;
  wire \nand_7.in_0 ;
  wire \nand_7.in_1 ;
  wire \nand_7.in_2 ;
  wire \nand_7.in_3 ;
  wire \nand_7.in_4 ;
  wire \nand_7.in_5 ;
  wire \nand_7.in_6 ;
  wire \nand_7.nand_0 ;
  wire \nand_7.nand_1 ;
  wire \nand_7.nand_2 ;
  wire \nand_7.nand_3 ;
  wire \nand_7.nand_4 ;
  wire \nand_7.out ;
  wire \nand_8.and_0 ;
  wire \nand_8.and_1 ;
  wire \nand_8.and_2 ;
  wire \nand_8.and_3 ;
  wire \nand_8.and_4 ;
  wire \nand_8.in_0 ;
  wire \nand_8.in_1 ;
  wire \nand_8.in_2 ;
  wire \nand_8.in_3 ;
  wire \nand_8.in_4 ;
  wire \nand_8.in_5 ;
  wire \nand_8.in_6 ;
  wire \nand_8.nand_0 ;
  wire \nand_8.nand_1 ;
  wire \nand_8.nand_2 ;
  wire \nand_8.nand_3 ;
  wire \nand_8.nand_4 ;
  wire \nand_8.out ;
  wire \nand_9.and_0 ;
  wire \nand_9.and_1 ;
  wire \nand_9.and_2 ;
  wire \nand_9.and_3 ;
  wire \nand_9.and_4 ;
  wire \nand_9.in_0 ;
  wire \nand_9.in_1 ;
  wire \nand_9.in_2 ;
  wire \nand_9.in_3 ;
  wire \nand_9.in_4 ;
  wire \nand_9.in_5 ;
  wire \nand_9.in_6 ;
  wire \nand_9.nand_0 ;
  wire \nand_9.nand_1 ;
  wire \nand_9.nand_2 ;
  wire \nand_9.nand_3 ;
  wire \nand_9.nand_4 ;
  wire \nand_9.out ;
  output \out<0> ;
  output \out<10> ;
  output \out<11> ;
  output \out<12> ;
  output \out<13> ;
  output \out<14> ;
  output \out<15> ;
  output \out<16> ;
  output \out<17> ;
  output \out<18> ;
  output \out<19> ;
  output \out<1> ;
  output \out<20> ;
  output \out<21> ;
  output \out<22> ;
  output \out<23> ;
  output \out<24> ;
  output \out<25> ;
  output \out<26> ;
  output \out<27> ;
  output \out<28> ;
  output \out<29> ;
  output \out<2> ;
  output \out<30> ;
  output \out<31> ;
  output \out<32> ;
  output \out<33> ;
  output \out<34> ;
  output \out<35> ;
  output \out<36> ;
  output \out<37> ;
  output \out<38> ;
  output \out<39> ;
  output \out<3> ;
  output \out<40> ;
  output \out<41> ;
  output \out<42> ;
  output \out<43> ;
  output \out<44> ;
  output \out<45> ;
  output \out<46> ;
  output \out<47> ;
  output \out<48> ;
  output \out<49> ;
  output \out<4> ;
  output \out<50> ;
  output \out<51> ;
  output \out<52> ;
  output \out<53> ;
  output \out<54> ;
  output \out<55> ;
  output \out<56> ;
  output \out<57> ;
  output \out<58> ;
  output \out<59> ;
  output \out<5> ;
  output \out<60> ;
  output \out<61> ;
  output \out<62> ;
  output \out<63> ;
  output \out<6> ;
  output \out<7> ;
  output \out<8> ;
  output \out<9> ;
  wire \out_b<0> ;
  wire \out_b<10> ;
  wire \out_b<11> ;
  wire \out_b<12> ;
  wire \out_b<13> ;
  wire \out_b<14> ;
  wire \out_b<15> ;
  wire \out_b<16> ;
  wire \out_b<17> ;
  wire \out_b<18> ;
  wire \out_b<19> ;
  wire \out_b<1> ;
  wire \out_b<20> ;
  wire \out_b<21> ;
  wire \out_b<22> ;
  wire \out_b<23> ;
  wire \out_b<24> ;
  wire \out_b<25> ;
  wire \out_b<26> ;
  wire \out_b<27> ;
  wire \out_b<28> ;
  wire \out_b<29> ;
  wire \out_b<2> ;
  wire \out_b<30> ;
  wire \out_b<31> ;
  wire \out_b<32> ;
  wire \out_b<33> ;
  wire \out_b<34> ;
  wire \out_b<35> ;
  wire \out_b<36> ;
  wire \out_b<37> ;
  wire \out_b<38> ;
  wire \out_b<39> ;
  wire \out_b<3> ;
  wire \out_b<40> ;
  wire \out_b<41> ;
  wire \out_b<42> ;
  wire \out_b<43> ;
  wire \out_b<44> ;
  wire \out_b<45> ;
  wire \out_b<46> ;
  wire \out_b<47> ;
  wire \out_b<48> ;
  wire \out_b<49> ;
  wire \out_b<4> ;
  wire \out_b<50> ;
  wire \out_b<51> ;
  wire \out_b<52> ;
  wire \out_b<53> ;
  wire \out_b<54> ;
  wire \out_b<55> ;
  wire \out_b<56> ;
  wire \out_b<57> ;
  wire \out_b<58> ;
  wire \out_b<59> ;
  wire \out_b<5> ;
  wire \out_b<60> ;
  wire \out_b<61> ;
  wire \out_b<62> ;
  wire \out_b<63> ;
  wire \out_b<6> ;
  wire \out_b<7> ;
  wire \out_b<8> ;
  wire \out_b<9> ;
  inverter inv_for_input_0 (    .in(\in<0> ),    .out(\in_b<0> )
  );
  inverter inv_for_input_1 (    .in(\in<1> ),    .out(\in_b<1> )
  );
  inverter inv_for_input_2 (    .in(\in<2> ),    .out(\in_b<2> )
  );
  inverter inv_for_input_3 (    .in(\in<3> ),    .out(\in_b<3> )
  );
  inverter inv_for_input_4 (    .in(\in<4> ),    .out(\in_b<4> )
  );
  inverter inv_for_input_5 (    .in(\in<5> ),    .out(\in_b<5> )
  );
  inverter inv_for_output_0 (    .in(\nand_0.out ),    .out(\out<0> )
  );
  inverter inv_for_output_1 (    .in(\nand_1.out ),    .out(\out<1> )
  );
  inverter inv_for_output_10 (    .in(\nand_10.out ),    .out(\out<10> )
  );
  inverter inv_for_output_11 (    .in(\nand_11.out ),    .out(\out<11> )
  );
  inverter inv_for_output_12 (    .in(\nand_12.out ),    .out(\out<12> )
  );
  inverter inv_for_output_13 (    .in(\nand_13.out ),    .out(\out<13> )
  );
  inverter inv_for_output_14 (    .in(\nand_14.out ),    .out(\out<14> )
  );
  inverter inv_for_output_15 (    .in(\nand_15.out ),    .out(\out<15> )
  );
  inverter inv_for_output_16 (    .in(\nand_16.out ),    .out(\out<16> )
  );
  inverter inv_for_output_17 (    .in(\nand_17.out ),    .out(\out<17> )
  );
  inverter inv_for_output_18 (    .in(\nand_18.out ),    .out(\out<18> )
  );
  inverter inv_for_output_19 (    .in(\nand_19.out ),    .out(\out<19> )
  );
  inverter inv_for_output_2 (    .in(\nand_2.out ),    .out(\out<2> )
  );
  inverter inv_for_output_20 (    .in(\nand_20.out ),    .out(\out<20> )
  );
  inverter inv_for_output_21 (    .in(\nand_21.out ),    .out(\out<21> )
  );
  inverter inv_for_output_22 (    .in(\nand_22.out ),    .out(\out<22> )
  );
  inverter inv_for_output_23 (    .in(\nand_23.out ),    .out(\out<23> )
  );
  inverter inv_for_output_24 (    .in(\nand_24.out ),    .out(\out<24> )
  );
  inverter inv_for_output_25 (    .in(\nand_25.out ),    .out(\out<25> )
  );
  inverter inv_for_output_26 (    .in(\nand_26.out ),    .out(\out<26> )
  );
  inverter inv_for_output_27 (    .in(\nand_27.out ),    .out(\out<27> )
  );
  inverter inv_for_output_28 (    .in(\nand_28.out ),    .out(\out<28> )
  );
  inverter inv_for_output_29 (    .in(\nand_29.out ),    .out(\out<29> )
  );
  inverter inv_for_output_3 (    .in(\nand_3.out ),    .out(\out<3> )
  );
  inverter inv_for_output_30 (    .in(\nand_30.out ),    .out(\out<30> )
  );
  inverter inv_for_output_31 (    .in(\nand_31.out ),    .out(\out<31> )
  );
  inverter inv_for_output_32 (    .in(\nand_32.out ),    .out(\out<32> )
  );
  inverter inv_for_output_33 (    .in(\nand_33.out ),    .out(\out<33> )
  );
  inverter inv_for_output_34 (    .in(\nand_34.out ),    .out(\out<34> )
  );
  inverter inv_for_output_35 (    .in(\nand_35.out ),    .out(\out<35> )
  );
  inverter inv_for_output_36 (    .in(\nand_36.out ),    .out(\out<36> )
  );
  inverter inv_for_output_37 (    .in(\nand_37.out ),    .out(\out<37> )
  );
  inverter inv_for_output_38 (    .in(\nand_38.out ),    .out(\out<38> )
  );
  inverter inv_for_output_39 (    .in(\nand_39.out ),    .out(\out<39> )
  );
  inverter inv_for_output_4 (    .in(\nand_4.out ),    .out(\out<4> )
  );
  inverter inv_for_output_40 (    .in(\nand_40.out ),    .out(\out<40> )
  );
  inverter inv_for_output_41 (    .in(\nand_41.out ),    .out(\out<41> )
  );
  inverter inv_for_output_42 (    .in(\nand_42.out ),    .out(\out<42> )
  );
  inverter inv_for_output_43 (    .in(\nand_43.out ),    .out(\out<43> )
  );
  inverter inv_for_output_44 (    .in(\nand_44.out ),    .out(\out<44> )
  );
  inverter inv_for_output_45 (    .in(\nand_45.out ),    .out(\out<45> )
  );
  inverter inv_for_output_46 (    .in(\nand_46.out ),    .out(\out<46> )
  );
  inverter inv_for_output_47 (    .in(\nand_47.out ),    .out(\out<47> )
  );
  inverter inv_for_output_48 (    .in(\nand_48.out ),    .out(\out<48> )
  );
  inverter inv_for_output_49 (    .in(\nand_49.out ),    .out(\out<49> )
  );
  inverter inv_for_output_5 (    .in(\nand_5.out ),    .out(\out<5> )
  );
  inverter inv_for_output_50 (    .in(\nand_50.out ),    .out(\out<50> )
  );
  inverter inv_for_output_51 (    .in(\nand_51.out ),    .out(\out<51> )
  );
  inverter inv_for_output_52 (    .in(\nand_52.out ),    .out(\out<52> )
  );
  inverter inv_for_output_53 (    .in(\nand_53.out ),    .out(\out<53> )
  );
  inverter inv_for_output_54 (    .in(\nand_54.out ),    .out(\out<54> )
  );
  inverter inv_for_output_55 (    .in(\nand_55.out ),    .out(\out<55> )
  );
  inverter inv_for_output_56 (    .in(\nand_56.out ),    .out(\out<56> )
  );
  inverter inv_for_output_57 (    .in(\nand_57.out ),    .out(\out<57> )
  );
  inverter inv_for_output_58 (    .in(\nand_58.out ),    .out(\out<58> )
  );
  inverter inv_for_output_59 (    .in(\nand_59.out ),    .out(\out<59> )
  );
  inverter inv_for_output_6 (    .in(\nand_6.out ),    .out(\out<6> )
  );
  inverter inv_for_output_60 (    .in(\nand_60.out ),    .out(\out<60> )
  );
  inverter inv_for_output_61 (    .in(\nand_61.out ),    .out(\out<61> )
  );
  inverter inv_for_output_62 (    .in(\nand_62.out ),    .out(\out<62> )
  );
  inverter inv_for_output_63 (    .in(\nand_63.out ),    .out(\out<63> )
  );
  inverter inv_for_output_7 (    .in(\nand_7.out ),    .out(\out<7> )
  );
  inverter inv_for_output_8 (    .in(\nand_8.out ),    .out(\out<8> )
  );
  inverter inv_for_output_9 (    .in(\nand_9.out ),    .out(\out<9> )
  );
  inverter \nand_0.inv_0  (    .in(\nand_0.nand_0 ),    .out(\nand_0.and_0 )
  );
  inverter \nand_0.inv_1  (    .in(\nand_0.nand_1 ),    .out(\nand_0.and_1 )
  );
  inverter \nand_0.inv_2  (    .in(\nand_0.nand_2 ),    .out(\nand_0.and_2 )
  );
  inverter \nand_0.inv_3  (    .in(\nand_0.nand_3 ),    .out(\nand_0.and_3 )
  );
  inverter \nand_0.inv_4  (    .in(\nand_0.nand_4 ),    .out(\nand_0.and_4 )
  );
  nand2 \nand_0.nand2_0  (    .in_0(\in_b<0> ),    .in_1(\in_b<1> ),    .out(\nand_0.nand_0 )
  );
  nand2 \nand_0.nand2_1  (    .in_0(\nand_0.and_0 ),    .in_1(\in_b<2> ),    .out(\nand_0.nand_1 )
  );
  nand2 \nand_0.nand2_2  (    .in_0(\nand_0.and_1 ),    .in_1(\in_b<3> ),    .out(\nand_0.nand_2 )
  );
  nand2 \nand_0.nand2_3  (    .in_0(\nand_0.and_2 ),    .in_1(\in_b<4> ),    .out(\nand_0.nand_3 )
  );
  nand2 \nand_0.nand2_4  (    .in_0(\nand_0.and_3 ),    .in_1(\in_b<5> ),    .out(\nand_0.nand_4 )
  );
  nand2 \nand_0.nand2_5  (    .in_0(\nand_0.and_4 ),    .in_1(enable),    .out(\nand_0.out )
  );
  inverter \nand_1.inv_0  (    .in(\nand_1.nand_0 ),    .out(\nand_1.and_0 )
  );
  inverter \nand_1.inv_1  (    .in(\nand_1.nand_1 ),    .out(\nand_1.and_1 )
  );
  inverter \nand_1.inv_2  (    .in(\nand_1.nand_2 ),    .out(\nand_1.and_2 )
  );
  inverter \nand_1.inv_3  (    .in(\nand_1.nand_3 ),    .out(\nand_1.and_3 )
  );
  inverter \nand_1.inv_4  (    .in(\nand_1.nand_4 ),    .out(\nand_1.and_4 )
  );
  nand2 \nand_1.nand2_0  (    .in_0(\in<0> ),    .in_1(\in_b<1> ),    .out(\nand_1.nand_0 )
  );
  nand2 \nand_1.nand2_1  (    .in_0(\nand_1.and_0 ),    .in_1(\in_b<2> ),    .out(\nand_1.nand_1 )
  );
  nand2 \nand_1.nand2_2  (    .in_0(\nand_1.and_1 ),    .in_1(\in_b<3> ),    .out(\nand_1.nand_2 )
  );
  nand2 \nand_1.nand2_3  (    .in_0(\nand_1.and_2 ),    .in_1(\in_b<4> ),    .out(\nand_1.nand_3 )
  );
  nand2 \nand_1.nand2_4  (    .in_0(\nand_1.and_3 ),    .in_1(\in_b<5> ),    .out(\nand_1.nand_4 )
  );
  nand2 \nand_1.nand2_5  (    .in_0(\nand_1.and_4 ),    .in_1(enable),    .out(\nand_1.out )
  );
  inverter \nand_10.inv_0  (    .in(\nand_10.nand_0 ),    .out(\nand_10.and_0 )
  );
  inverter \nand_10.inv_1  (    .in(\nand_10.nand_1 ),    .out(\nand_10.and_1 )
  );
  inverter \nand_10.inv_2  (    .in(\nand_10.nand_2 ),    .out(\nand_10.and_2 )
  );
  inverter \nand_10.inv_3  (    .in(\nand_10.nand_3 ),    .out(\nand_10.and_3 )
  );
  inverter \nand_10.inv_4  (    .in(\nand_10.nand_4 ),    .out(\nand_10.and_4 )
  );
  nand2 \nand_10.nand2_0  (    .in_0(\in_b<0> ),    .in_1(\in<1> ),    .out(\nand_10.nand_0 )
  );
  nand2 \nand_10.nand2_1  (    .in_0(\nand_10.and_0 ),    .in_1(\in_b<2> ),    .out(\nand_10.nand_1 )
  );
  nand2 \nand_10.nand2_2  (    .in_0(\nand_10.and_1 ),    .in_1(\in<3> ),    .out(\nand_10.nand_2 )
  );
  nand2 \nand_10.nand2_3  (    .in_0(\nand_10.and_2 ),    .in_1(\in_b<4> ),    .out(\nand_10.nand_3 )
  );
  nand2 \nand_10.nand2_4  (    .in_0(\nand_10.and_3 ),    .in_1(\in_b<5> ),    .out(\nand_10.nand_4 )
  );
  nand2 \nand_10.nand2_5  (    .in_0(\nand_10.and_4 ),    .in_1(enable),    .out(\nand_10.out )
  );
  inverter \nand_11.inv_0  (    .in(\nand_11.nand_0 ),    .out(\nand_11.and_0 )
  );
  inverter \nand_11.inv_1  (    .in(\nand_11.nand_1 ),    .out(\nand_11.and_1 )
  );
  inverter \nand_11.inv_2  (    .in(\nand_11.nand_2 ),    .out(\nand_11.and_2 )
  );
  inverter \nand_11.inv_3  (    .in(\nand_11.nand_3 ),    .out(\nand_11.and_3 )
  );
  inverter \nand_11.inv_4  (    .in(\nand_11.nand_4 ),    .out(\nand_11.and_4 )
  );
  nand2 \nand_11.nand2_0  (    .in_0(\in<0> ),    .in_1(\in<1> ),    .out(\nand_11.nand_0 )
  );
  nand2 \nand_11.nand2_1  (    .in_0(\nand_11.and_0 ),    .in_1(\in_b<2> ),    .out(\nand_11.nand_1 )
  );
  nand2 \nand_11.nand2_2  (    .in_0(\nand_11.and_1 ),    .in_1(\in<3> ),    .out(\nand_11.nand_2 )
  );
  nand2 \nand_11.nand2_3  (    .in_0(\nand_11.and_2 ),    .in_1(\in_b<4> ),    .out(\nand_11.nand_3 )
  );
  nand2 \nand_11.nand2_4  (    .in_0(\nand_11.and_3 ),    .in_1(\in_b<5> ),    .out(\nand_11.nand_4 )
  );
  nand2 \nand_11.nand2_5  (    .in_0(\nand_11.and_4 ),    .in_1(enable),    .out(\nand_11.out )
  );
  inverter \nand_12.inv_0  (    .in(\nand_12.nand_0 ),    .out(\nand_12.and_0 )
  );
  inverter \nand_12.inv_1  (    .in(\nand_12.nand_1 ),    .out(\nand_12.and_1 )
  );
  inverter \nand_12.inv_2  (    .in(\nand_12.nand_2 ),    .out(\nand_12.and_2 )
  );
  inverter \nand_12.inv_3  (    .in(\nand_12.nand_3 ),    .out(\nand_12.and_3 )
  );
  inverter \nand_12.inv_4  (    .in(\nand_12.nand_4 ),    .out(\nand_12.and_4 )
  );
  nand2 \nand_12.nand2_0  (    .in_0(\in_b<0> ),    .in_1(\in_b<1> ),    .out(\nand_12.nand_0 )
  );
  nand2 \nand_12.nand2_1  (    .in_0(\nand_12.and_0 ),    .in_1(\in<2> ),    .out(\nand_12.nand_1 )
  );
  nand2 \nand_12.nand2_2  (    .in_0(\nand_12.and_1 ),    .in_1(\in<3> ),    .out(\nand_12.nand_2 )
  );
  nand2 \nand_12.nand2_3  (    .in_0(\nand_12.and_2 ),    .in_1(\in_b<4> ),    .out(\nand_12.nand_3 )
  );
  nand2 \nand_12.nand2_4  (    .in_0(\nand_12.and_3 ),    .in_1(\in_b<5> ),    .out(\nand_12.nand_4 )
  );
  nand2 \nand_12.nand2_5  (    .in_0(\nand_12.and_4 ),    .in_1(enable),    .out(\nand_12.out )
  );
  inverter \nand_13.inv_0  (    .in(\nand_13.nand_0 ),    .out(\nand_13.and_0 )
  );
  inverter \nand_13.inv_1  (    .in(\nand_13.nand_1 ),    .out(\nand_13.and_1 )
  );
  inverter \nand_13.inv_2  (    .in(\nand_13.nand_2 ),    .out(\nand_13.and_2 )
  );
  inverter \nand_13.inv_3  (    .in(\nand_13.nand_3 ),    .out(\nand_13.and_3 )
  );
  inverter \nand_13.inv_4  (    .in(\nand_13.nand_4 ),    .out(\nand_13.and_4 )
  );
  nand2 \nand_13.nand2_0  (    .in_0(\in<0> ),    .in_1(\in_b<1> ),    .out(\nand_13.nand_0 )
  );
  nand2 \nand_13.nand2_1  (    .in_0(\nand_13.and_0 ),    .in_1(\in<2> ),    .out(\nand_13.nand_1 )
  );
  nand2 \nand_13.nand2_2  (    .in_0(\nand_13.and_1 ),    .in_1(\in<3> ),    .out(\nand_13.nand_2 )
  );
  nand2 \nand_13.nand2_3  (    .in_0(\nand_13.and_2 ),    .in_1(\in_b<4> ),    .out(\nand_13.nand_3 )
  );
  nand2 \nand_13.nand2_4  (    .in_0(\nand_13.and_3 ),    .in_1(\in_b<5> ),    .out(\nand_13.nand_4 )
  );
  nand2 \nand_13.nand2_5  (    .in_0(\nand_13.and_4 ),    .in_1(enable),    .out(\nand_13.out )
  );
  inverter \nand_14.inv_0  (    .in(\nand_14.nand_0 ),    .out(\nand_14.and_0 )
  );
  inverter \nand_14.inv_1  (    .in(\nand_14.nand_1 ),    .out(\nand_14.and_1 )
  );
  inverter \nand_14.inv_2  (    .in(\nand_14.nand_2 ),    .out(\nand_14.and_2 )
  );
  inverter \nand_14.inv_3  (    .in(\nand_14.nand_3 ),    .out(\nand_14.and_3 )
  );
  inverter \nand_14.inv_4  (    .in(\nand_14.nand_4 ),    .out(\nand_14.and_4 )
  );
  nand2 \nand_14.nand2_0  (    .in_0(\in_b<0> ),    .in_1(\in<1> ),    .out(\nand_14.nand_0 )
  );
  nand2 \nand_14.nand2_1  (    .in_0(\nand_14.and_0 ),    .in_1(\in<2> ),    .out(\nand_14.nand_1 )
  );
  nand2 \nand_14.nand2_2  (    .in_0(\nand_14.and_1 ),    .in_1(\in<3> ),    .out(\nand_14.nand_2 )
  );
  nand2 \nand_14.nand2_3  (    .in_0(\nand_14.and_2 ),    .in_1(\in_b<4> ),    .out(\nand_14.nand_3 )
  );
  nand2 \nand_14.nand2_4  (    .in_0(\nand_14.and_3 ),    .in_1(\in_b<5> ),    .out(\nand_14.nand_4 )
  );
  nand2 \nand_14.nand2_5  (    .in_0(\nand_14.and_4 ),    .in_1(enable),    .out(\nand_14.out )
  );
  inverter \nand_15.inv_0  (    .in(\nand_15.nand_0 ),    .out(\nand_15.and_0 )
  );
  inverter \nand_15.inv_1  (    .in(\nand_15.nand_1 ),    .out(\nand_15.and_1 )
  );
  inverter \nand_15.inv_2  (    .in(\nand_15.nand_2 ),    .out(\nand_15.and_2 )
  );
  inverter \nand_15.inv_3  (    .in(\nand_15.nand_3 ),    .out(\nand_15.and_3 )
  );
  inverter \nand_15.inv_4  (    .in(\nand_15.nand_4 ),    .out(\nand_15.and_4 )
  );
  nand2 \nand_15.nand2_0  (    .in_0(\in<0> ),    .in_1(\in<1> ),    .out(\nand_15.nand_0 )
  );
  nand2 \nand_15.nand2_1  (    .in_0(\nand_15.and_0 ),    .in_1(\in<2> ),    .out(\nand_15.nand_1 )
  );
  nand2 \nand_15.nand2_2  (    .in_0(\nand_15.and_1 ),    .in_1(\in<3> ),    .out(\nand_15.nand_2 )
  );
  nand2 \nand_15.nand2_3  (    .in_0(\nand_15.and_2 ),    .in_1(\in_b<4> ),    .out(\nand_15.nand_3 )
  );
  nand2 \nand_15.nand2_4  (    .in_0(\nand_15.and_3 ),    .in_1(\in_b<5> ),    .out(\nand_15.nand_4 )
  );
  nand2 \nand_15.nand2_5  (    .in_0(\nand_15.and_4 ),    .in_1(enable),    .out(\nand_15.out )
  );
  inverter \nand_16.inv_0  (    .in(\nand_16.nand_0 ),    .out(\nand_16.and_0 )
  );
  inverter \nand_16.inv_1  (    .in(\nand_16.nand_1 ),    .out(\nand_16.and_1 )
  );
  inverter \nand_16.inv_2  (    .in(\nand_16.nand_2 ),    .out(\nand_16.and_2 )
  );
  inverter \nand_16.inv_3  (    .in(\nand_16.nand_3 ),    .out(\nand_16.and_3 )
  );
  inverter \nand_16.inv_4  (    .in(\nand_16.nand_4 ),    .out(\nand_16.and_4 )
  );
  nand2 \nand_16.nand2_0  (    .in_0(\in_b<0> ),    .in_1(\in_b<1> ),    .out(\nand_16.nand_0 )
  );
  nand2 \nand_16.nand2_1  (    .in_0(\nand_16.and_0 ),    .in_1(\in_b<2> ),    .out(\nand_16.nand_1 )
  );
  nand2 \nand_16.nand2_2  (    .in_0(\nand_16.and_1 ),    .in_1(\in_b<3> ),    .out(\nand_16.nand_2 )
  );
  nand2 \nand_16.nand2_3  (    .in_0(\nand_16.and_2 ),    .in_1(\in<4> ),    .out(\nand_16.nand_3 )
  );
  nand2 \nand_16.nand2_4  (    .in_0(\nand_16.and_3 ),    .in_1(\in_b<5> ),    .out(\nand_16.nand_4 )
  );
  nand2 \nand_16.nand2_5  (    .in_0(\nand_16.and_4 ),    .in_1(enable),    .out(\nand_16.out )
  );
  inverter \nand_17.inv_0  (    .in(\nand_17.nand_0 ),    .out(\nand_17.and_0 )
  );
  inverter \nand_17.inv_1  (    .in(\nand_17.nand_1 ),    .out(\nand_17.and_1 )
  );
  inverter \nand_17.inv_2  (    .in(\nand_17.nand_2 ),    .out(\nand_17.and_2 )
  );
  inverter \nand_17.inv_3  (    .in(\nand_17.nand_3 ),    .out(\nand_17.and_3 )
  );
  inverter \nand_17.inv_4  (    .in(\nand_17.nand_4 ),    .out(\nand_17.and_4 )
  );
  nand2 \nand_17.nand2_0  (    .in_0(\in<0> ),    .in_1(\in_b<1> ),    .out(\nand_17.nand_0 )
  );
  nand2 \nand_17.nand2_1  (    .in_0(\nand_17.and_0 ),    .in_1(\in_b<2> ),    .out(\nand_17.nand_1 )
  );
  nand2 \nand_17.nand2_2  (    .in_0(\nand_17.and_1 ),    .in_1(\in_b<3> ),    .out(\nand_17.nand_2 )
  );
  nand2 \nand_17.nand2_3  (    .in_0(\nand_17.and_2 ),    .in_1(\in<4> ),    .out(\nand_17.nand_3 )
  );
  nand2 \nand_17.nand2_4  (    .in_0(\nand_17.and_3 ),    .in_1(\in_b<5> ),    .out(\nand_17.nand_4 )
  );
  nand2 \nand_17.nand2_5  (    .in_0(\nand_17.and_4 ),    .in_1(enable),    .out(\nand_17.out )
  );
  inverter \nand_18.inv_0  (    .in(\nand_18.nand_0 ),    .out(\nand_18.and_0 )
  );
  inverter \nand_18.inv_1  (    .in(\nand_18.nand_1 ),    .out(\nand_18.and_1 )
  );
  inverter \nand_18.inv_2  (    .in(\nand_18.nand_2 ),    .out(\nand_18.and_2 )
  );
  inverter \nand_18.inv_3  (    .in(\nand_18.nand_3 ),    .out(\nand_18.and_3 )
  );
  inverter \nand_18.inv_4  (    .in(\nand_18.nand_4 ),    .out(\nand_18.and_4 )
  );
  nand2 \nand_18.nand2_0  (    .in_0(\in_b<0> ),    .in_1(\in<1> ),    .out(\nand_18.nand_0 )
  );
  nand2 \nand_18.nand2_1  (    .in_0(\nand_18.and_0 ),    .in_1(\in_b<2> ),    .out(\nand_18.nand_1 )
  );
  nand2 \nand_18.nand2_2  (    .in_0(\nand_18.and_1 ),    .in_1(\in_b<3> ),    .out(\nand_18.nand_2 )
  );
  nand2 \nand_18.nand2_3  (    .in_0(\nand_18.and_2 ),    .in_1(\in<4> ),    .out(\nand_18.nand_3 )
  );
  nand2 \nand_18.nand2_4  (    .in_0(\nand_18.and_3 ),    .in_1(\in_b<5> ),    .out(\nand_18.nand_4 )
  );
  nand2 \nand_18.nand2_5  (    .in_0(\nand_18.and_4 ),    .in_1(enable),    .out(\nand_18.out )
  );
  inverter \nand_19.inv_0  (    .in(\nand_19.nand_0 ),    .out(\nand_19.and_0 )
  );
  inverter \nand_19.inv_1  (    .in(\nand_19.nand_1 ),    .out(\nand_19.and_1 )
  );
  inverter \nand_19.inv_2  (    .in(\nand_19.nand_2 ),    .out(\nand_19.and_2 )
  );
  inverter \nand_19.inv_3  (    .in(\nand_19.nand_3 ),    .out(\nand_19.and_3 )
  );
  inverter \nand_19.inv_4  (    .in(\nand_19.nand_4 ),    .out(\nand_19.and_4 )
  );
  nand2 \nand_19.nand2_0  (    .in_0(\in<0> ),    .in_1(\in<1> ),    .out(\nand_19.nand_0 )
  );
  nand2 \nand_19.nand2_1  (    .in_0(\nand_19.and_0 ),    .in_1(\in_b<2> ),    .out(\nand_19.nand_1 )
  );
  nand2 \nand_19.nand2_2  (    .in_0(\nand_19.and_1 ),    .in_1(\in_b<3> ),    .out(\nand_19.nand_2 )
  );
  nand2 \nand_19.nand2_3  (    .in_0(\nand_19.and_2 ),    .in_1(\in<4> ),    .out(\nand_19.nand_3 )
  );
  nand2 \nand_19.nand2_4  (    .in_0(\nand_19.and_3 ),    .in_1(\in_b<5> ),    .out(\nand_19.nand_4 )
  );
  nand2 \nand_19.nand2_5  (    .in_0(\nand_19.and_4 ),    .in_1(enable),    .out(\nand_19.out )
  );
  inverter \nand_2.inv_0  (    .in(\nand_2.nand_0 ),    .out(\nand_2.and_0 )
  );
  inverter \nand_2.inv_1  (    .in(\nand_2.nand_1 ),    .out(\nand_2.and_1 )
  );
  inverter \nand_2.inv_2  (    .in(\nand_2.nand_2 ),    .out(\nand_2.and_2 )
  );
  inverter \nand_2.inv_3  (    .in(\nand_2.nand_3 ),    .out(\nand_2.and_3 )
  );
  inverter \nand_2.inv_4  (    .in(\nand_2.nand_4 ),    .out(\nand_2.and_4 )
  );
  nand2 \nand_2.nand2_0  (    .in_0(\in_b<0> ),    .in_1(\in<1> ),    .out(\nand_2.nand_0 )
  );
  nand2 \nand_2.nand2_1  (    .in_0(\nand_2.and_0 ),    .in_1(\in_b<2> ),    .out(\nand_2.nand_1 )
  );
  nand2 \nand_2.nand2_2  (    .in_0(\nand_2.and_1 ),    .in_1(\in_b<3> ),    .out(\nand_2.nand_2 )
  );
  nand2 \nand_2.nand2_3  (    .in_0(\nand_2.and_2 ),    .in_1(\in_b<4> ),    .out(\nand_2.nand_3 )
  );
  nand2 \nand_2.nand2_4  (    .in_0(\nand_2.and_3 ),    .in_1(\in_b<5> ),    .out(\nand_2.nand_4 )
  );
  nand2 \nand_2.nand2_5  (    .in_0(\nand_2.and_4 ),    .in_1(enable),    .out(\nand_2.out )
  );
  inverter \nand_20.inv_0  (    .in(\nand_20.nand_0 ),    .out(\nand_20.and_0 )
  );
  inverter \nand_20.inv_1  (    .in(\nand_20.nand_1 ),    .out(\nand_20.and_1 )
  );
  inverter \nand_20.inv_2  (    .in(\nand_20.nand_2 ),    .out(\nand_20.and_2 )
  );
  inverter \nand_20.inv_3  (    .in(\nand_20.nand_3 ),    .out(\nand_20.and_3 )
  );
  inverter \nand_20.inv_4  (    .in(\nand_20.nand_4 ),    .out(\nand_20.and_4 )
  );
  nand2 \nand_20.nand2_0  (    .in_0(\in_b<0> ),    .in_1(\in_b<1> ),    .out(\nand_20.nand_0 )
  );
  nand2 \nand_20.nand2_1  (    .in_0(\nand_20.and_0 ),    .in_1(\in<2> ),    .out(\nand_20.nand_1 )
  );
  nand2 \nand_20.nand2_2  (    .in_0(\nand_20.and_1 ),    .in_1(\in_b<3> ),    .out(\nand_20.nand_2 )
  );
  nand2 \nand_20.nand2_3  (    .in_0(\nand_20.and_2 ),    .in_1(\in<4> ),    .out(\nand_20.nand_3 )
  );
  nand2 \nand_20.nand2_4  (    .in_0(\nand_20.and_3 ),    .in_1(\in_b<5> ),    .out(\nand_20.nand_4 )
  );
  nand2 \nand_20.nand2_5  (    .in_0(\nand_20.and_4 ),    .in_1(enable),    .out(\nand_20.out )
  );
  inverter \nand_21.inv_0  (    .in(\nand_21.nand_0 ),    .out(\nand_21.and_0 )
  );
  inverter \nand_21.inv_1  (    .in(\nand_21.nand_1 ),    .out(\nand_21.and_1 )
  );
  inverter \nand_21.inv_2  (    .in(\nand_21.nand_2 ),    .out(\nand_21.and_2 )
  );
  inverter \nand_21.inv_3  (    .in(\nand_21.nand_3 ),    .out(\nand_21.and_3 )
  );
  inverter \nand_21.inv_4  (    .in(\nand_21.nand_4 ),    .out(\nand_21.and_4 )
  );
  nand2 \nand_21.nand2_0  (    .in_0(\in<0> ),    .in_1(\in_b<1> ),    .out(\nand_21.nand_0 )
  );
  nand2 \nand_21.nand2_1  (    .in_0(\nand_21.and_0 ),    .in_1(\in<2> ),    .out(\nand_21.nand_1 )
  );
  nand2 \nand_21.nand2_2  (    .in_0(\nand_21.and_1 ),    .in_1(\in_b<3> ),    .out(\nand_21.nand_2 )
  );
  nand2 \nand_21.nand2_3  (    .in_0(\nand_21.and_2 ),    .in_1(\in<4> ),    .out(\nand_21.nand_3 )
  );
  nand2 \nand_21.nand2_4  (    .in_0(\nand_21.and_3 ),    .in_1(\in_b<5> ),    .out(\nand_21.nand_4 )
  );
  nand2 \nand_21.nand2_5  (    .in_0(\nand_21.and_4 ),    .in_1(enable),    .out(\nand_21.out )
  );
  inverter \nand_22.inv_0  (    .in(\nand_22.nand_0 ),    .out(\nand_22.and_0 )
  );
  inverter \nand_22.inv_1  (    .in(\nand_22.nand_1 ),    .out(\nand_22.and_1 )
  );
  inverter \nand_22.inv_2  (    .in(\nand_22.nand_2 ),    .out(\nand_22.and_2 )
  );
  inverter \nand_22.inv_3  (    .in(\nand_22.nand_3 ),    .out(\nand_22.and_3 )
  );
  inverter \nand_22.inv_4  (    .in(\nand_22.nand_4 ),    .out(\nand_22.and_4 )
  );
  nand2 \nand_22.nand2_0  (    .in_0(\in_b<0> ),    .in_1(\in<1> ),    .out(\nand_22.nand_0 )
  );
  nand2 \nand_22.nand2_1  (    .in_0(\nand_22.and_0 ),    .in_1(\in<2> ),    .out(\nand_22.nand_1 )
  );
  nand2 \nand_22.nand2_2  (    .in_0(\nand_22.and_1 ),    .in_1(\in_b<3> ),    .out(\nand_22.nand_2 )
  );
  nand2 \nand_22.nand2_3  (    .in_0(\nand_22.and_2 ),    .in_1(\in<4> ),    .out(\nand_22.nand_3 )
  );
  nand2 \nand_22.nand2_4  (    .in_0(\nand_22.and_3 ),    .in_1(\in_b<5> ),    .out(\nand_22.nand_4 )
  );
  nand2 \nand_22.nand2_5  (    .in_0(\nand_22.and_4 ),    .in_1(enable),    .out(\nand_22.out )
  );
  inverter \nand_23.inv_0  (    .in(\nand_23.nand_0 ),    .out(\nand_23.and_0 )
  );
  inverter \nand_23.inv_1  (    .in(\nand_23.nand_1 ),    .out(\nand_23.and_1 )
  );
  inverter \nand_23.inv_2  (    .in(\nand_23.nand_2 ),    .out(\nand_23.and_2 )
  );
  inverter \nand_23.inv_3  (    .in(\nand_23.nand_3 ),    .out(\nand_23.and_3 )
  );
  inverter \nand_23.inv_4  (    .in(\nand_23.nand_4 ),    .out(\nand_23.and_4 )
  );
  nand2 \nand_23.nand2_0  (    .in_0(\in<0> ),    .in_1(\in<1> ),    .out(\nand_23.nand_0 )
  );
  nand2 \nand_23.nand2_1  (    .in_0(\nand_23.and_0 ),    .in_1(\in<2> ),    .out(\nand_23.nand_1 )
  );
  nand2 \nand_23.nand2_2  (    .in_0(\nand_23.and_1 ),    .in_1(\in_b<3> ),    .out(\nand_23.nand_2 )
  );
  nand2 \nand_23.nand2_3  (    .in_0(\nand_23.and_2 ),    .in_1(\in<4> ),    .out(\nand_23.nand_3 )
  );
  nand2 \nand_23.nand2_4  (    .in_0(\nand_23.and_3 ),    .in_1(\in_b<5> ),    .out(\nand_23.nand_4 )
  );
  nand2 \nand_23.nand2_5  (    .in_0(\nand_23.and_4 ),    .in_1(enable),    .out(\nand_23.out )
  );
  inverter \nand_24.inv_0  (    .in(\nand_24.nand_0 ),    .out(\nand_24.and_0 )
  );
  inverter \nand_24.inv_1  (    .in(\nand_24.nand_1 ),    .out(\nand_24.and_1 )
  );
  inverter \nand_24.inv_2  (    .in(\nand_24.nand_2 ),    .out(\nand_24.and_2 )
  );
  inverter \nand_24.inv_3  (    .in(\nand_24.nand_3 ),    .out(\nand_24.and_3 )
  );
  inverter \nand_24.inv_4  (    .in(\nand_24.nand_4 ),    .out(\nand_24.and_4 )
  );
  nand2 \nand_24.nand2_0  (    .in_0(\in_b<0> ),    .in_1(\in_b<1> ),    .out(\nand_24.nand_0 )
  );
  nand2 \nand_24.nand2_1  (    .in_0(\nand_24.and_0 ),    .in_1(\in_b<2> ),    .out(\nand_24.nand_1 )
  );
  nand2 \nand_24.nand2_2  (    .in_0(\nand_24.and_1 ),    .in_1(\in<3> ),    .out(\nand_24.nand_2 )
  );
  nand2 \nand_24.nand2_3  (    .in_0(\nand_24.and_2 ),    .in_1(\in<4> ),    .out(\nand_24.nand_3 )
  );
  nand2 \nand_24.nand2_4  (    .in_0(\nand_24.and_3 ),    .in_1(\in_b<5> ),    .out(\nand_24.nand_4 )
  );
  nand2 \nand_24.nand2_5  (    .in_0(\nand_24.and_4 ),    .in_1(enable),    .out(\nand_24.out )
  );
  inverter \nand_25.inv_0  (    .in(\nand_25.nand_0 ),    .out(\nand_25.and_0 )
  );
  inverter \nand_25.inv_1  (    .in(\nand_25.nand_1 ),    .out(\nand_25.and_1 )
  );
  inverter \nand_25.inv_2  (    .in(\nand_25.nand_2 ),    .out(\nand_25.and_2 )
  );
  inverter \nand_25.inv_3  (    .in(\nand_25.nand_3 ),    .out(\nand_25.and_3 )
  );
  inverter \nand_25.inv_4  (    .in(\nand_25.nand_4 ),    .out(\nand_25.and_4 )
  );
  nand2 \nand_25.nand2_0  (    .in_0(\in<0> ),    .in_1(\in_b<1> ),    .out(\nand_25.nand_0 )
  );
  nand2 \nand_25.nand2_1  (    .in_0(\nand_25.and_0 ),    .in_1(\in_b<2> ),    .out(\nand_25.nand_1 )
  );
  nand2 \nand_25.nand2_2  (    .in_0(\nand_25.and_1 ),    .in_1(\in<3> ),    .out(\nand_25.nand_2 )
  );
  nand2 \nand_25.nand2_3  (    .in_0(\nand_25.and_2 ),    .in_1(\in<4> ),    .out(\nand_25.nand_3 )
  );
  nand2 \nand_25.nand2_4  (    .in_0(\nand_25.and_3 ),    .in_1(\in_b<5> ),    .out(\nand_25.nand_4 )
  );
  nand2 \nand_25.nand2_5  (    .in_0(\nand_25.and_4 ),    .in_1(enable),    .out(\nand_25.out )
  );
  inverter \nand_26.inv_0  (    .in(\nand_26.nand_0 ),    .out(\nand_26.and_0 )
  );
  inverter \nand_26.inv_1  (    .in(\nand_26.nand_1 ),    .out(\nand_26.and_1 )
  );
  inverter \nand_26.inv_2  (    .in(\nand_26.nand_2 ),    .out(\nand_26.and_2 )
  );
  inverter \nand_26.inv_3  (    .in(\nand_26.nand_3 ),    .out(\nand_26.and_3 )
  );
  inverter \nand_26.inv_4  (    .in(\nand_26.nand_4 ),    .out(\nand_26.and_4 )
  );
  nand2 \nand_26.nand2_0  (    .in_0(\in_b<0> ),    .in_1(\in<1> ),    .out(\nand_26.nand_0 )
  );
  nand2 \nand_26.nand2_1  (    .in_0(\nand_26.and_0 ),    .in_1(\in_b<2> ),    .out(\nand_26.nand_1 )
  );
  nand2 \nand_26.nand2_2  (    .in_0(\nand_26.and_1 ),    .in_1(\in<3> ),    .out(\nand_26.nand_2 )
  );
  nand2 \nand_26.nand2_3  (    .in_0(\nand_26.and_2 ),    .in_1(\in<4> ),    .out(\nand_26.nand_3 )
  );
  nand2 \nand_26.nand2_4  (    .in_0(\nand_26.and_3 ),    .in_1(\in_b<5> ),    .out(\nand_26.nand_4 )
  );
  nand2 \nand_26.nand2_5  (    .in_0(\nand_26.and_4 ),    .in_1(enable),    .out(\nand_26.out )
  );
  inverter \nand_27.inv_0  (    .in(\nand_27.nand_0 ),    .out(\nand_27.and_0 )
  );
  inverter \nand_27.inv_1  (    .in(\nand_27.nand_1 ),    .out(\nand_27.and_1 )
  );
  inverter \nand_27.inv_2  (    .in(\nand_27.nand_2 ),    .out(\nand_27.and_2 )
  );
  inverter \nand_27.inv_3  (    .in(\nand_27.nand_3 ),    .out(\nand_27.and_3 )
  );
  inverter \nand_27.inv_4  (    .in(\nand_27.nand_4 ),    .out(\nand_27.and_4 )
  );
  nand2 \nand_27.nand2_0  (    .in_0(\in<0> ),    .in_1(\in<1> ),    .out(\nand_27.nand_0 )
  );
  nand2 \nand_27.nand2_1  (    .in_0(\nand_27.and_0 ),    .in_1(\in_b<2> ),    .out(\nand_27.nand_1 )
  );
  nand2 \nand_27.nand2_2  (    .in_0(\nand_27.and_1 ),    .in_1(\in<3> ),    .out(\nand_27.nand_2 )
  );
  nand2 \nand_27.nand2_3  (    .in_0(\nand_27.and_2 ),    .in_1(\in<4> ),    .out(\nand_27.nand_3 )
  );
  nand2 \nand_27.nand2_4  (    .in_0(\nand_27.and_3 ),    .in_1(\in_b<5> ),    .out(\nand_27.nand_4 )
  );
  nand2 \nand_27.nand2_5  (    .in_0(\nand_27.and_4 ),    .in_1(enable),    .out(\nand_27.out )
  );
  inverter \nand_28.inv_0  (    .in(\nand_28.nand_0 ),    .out(\nand_28.and_0 )
  );
  inverter \nand_28.inv_1  (    .in(\nand_28.nand_1 ),    .out(\nand_28.and_1 )
  );
  inverter \nand_28.inv_2  (    .in(\nand_28.nand_2 ),    .out(\nand_28.and_2 )
  );
  inverter \nand_28.inv_3  (    .in(\nand_28.nand_3 ),    .out(\nand_28.and_3 )
  );
  inverter \nand_28.inv_4  (    .in(\nand_28.nand_4 ),    .out(\nand_28.and_4 )
  );
  nand2 \nand_28.nand2_0  (    .in_0(\in_b<0> ),    .in_1(\in_b<1> ),    .out(\nand_28.nand_0 )
  );
  nand2 \nand_28.nand2_1  (    .in_0(\nand_28.and_0 ),    .in_1(\in<2> ),    .out(\nand_28.nand_1 )
  );
  nand2 \nand_28.nand2_2  (    .in_0(\nand_28.and_1 ),    .in_1(\in<3> ),    .out(\nand_28.nand_2 )
  );
  nand2 \nand_28.nand2_3  (    .in_0(\nand_28.and_2 ),    .in_1(\in<4> ),    .out(\nand_28.nand_3 )
  );
  nand2 \nand_28.nand2_4  (    .in_0(\nand_28.and_3 ),    .in_1(\in_b<5> ),    .out(\nand_28.nand_4 )
  );
  nand2 \nand_28.nand2_5  (    .in_0(\nand_28.and_4 ),    .in_1(enable),    .out(\nand_28.out )
  );
  inverter \nand_29.inv_0  (    .in(\nand_29.nand_0 ),    .out(\nand_29.and_0 )
  );
  inverter \nand_29.inv_1  (    .in(\nand_29.nand_1 ),    .out(\nand_29.and_1 )
  );
  inverter \nand_29.inv_2  (    .in(\nand_29.nand_2 ),    .out(\nand_29.and_2 )
  );
  inverter \nand_29.inv_3  (    .in(\nand_29.nand_3 ),    .out(\nand_29.and_3 )
  );
  inverter \nand_29.inv_4  (    .in(\nand_29.nand_4 ),    .out(\nand_29.and_4 )
  );
  nand2 \nand_29.nand2_0  (    .in_0(\in<0> ),    .in_1(\in_b<1> ),    .out(\nand_29.nand_0 )
  );
  nand2 \nand_29.nand2_1  (    .in_0(\nand_29.and_0 ),    .in_1(\in<2> ),    .out(\nand_29.nand_1 )
  );
  nand2 \nand_29.nand2_2  (    .in_0(\nand_29.and_1 ),    .in_1(\in<3> ),    .out(\nand_29.nand_2 )
  );
  nand2 \nand_29.nand2_3  (    .in_0(\nand_29.and_2 ),    .in_1(\in<4> ),    .out(\nand_29.nand_3 )
  );
  nand2 \nand_29.nand2_4  (    .in_0(\nand_29.and_3 ),    .in_1(\in_b<5> ),    .out(\nand_29.nand_4 )
  );
  nand2 \nand_29.nand2_5  (    .in_0(\nand_29.and_4 ),    .in_1(enable),    .out(\nand_29.out )
  );
  inverter \nand_3.inv_0  (    .in(\nand_3.nand_0 ),    .out(\nand_3.and_0 )
  );
  inverter \nand_3.inv_1  (    .in(\nand_3.nand_1 ),    .out(\nand_3.and_1 )
  );
  inverter \nand_3.inv_2  (    .in(\nand_3.nand_2 ),    .out(\nand_3.and_2 )
  );
  inverter \nand_3.inv_3  (    .in(\nand_3.nand_3 ),    .out(\nand_3.and_3 )
  );
  inverter \nand_3.inv_4  (    .in(\nand_3.nand_4 ),    .out(\nand_3.and_4 )
  );
  nand2 \nand_3.nand2_0  (    .in_0(\in<0> ),    .in_1(\in<1> ),    .out(\nand_3.nand_0 )
  );
  nand2 \nand_3.nand2_1  (    .in_0(\nand_3.and_0 ),    .in_1(\in_b<2> ),    .out(\nand_3.nand_1 )
  );
  nand2 \nand_3.nand2_2  (    .in_0(\nand_3.and_1 ),    .in_1(\in_b<3> ),    .out(\nand_3.nand_2 )
  );
  nand2 \nand_3.nand2_3  (    .in_0(\nand_3.and_2 ),    .in_1(\in_b<4> ),    .out(\nand_3.nand_3 )
  );
  nand2 \nand_3.nand2_4  (    .in_0(\nand_3.and_3 ),    .in_1(\in_b<5> ),    .out(\nand_3.nand_4 )
  );
  nand2 \nand_3.nand2_5  (    .in_0(\nand_3.and_4 ),    .in_1(enable),    .out(\nand_3.out )
  );
  inverter \nand_30.inv_0  (    .in(\nand_30.nand_0 ),    .out(\nand_30.and_0 )
  );
  inverter \nand_30.inv_1  (    .in(\nand_30.nand_1 ),    .out(\nand_30.and_1 )
  );
  inverter \nand_30.inv_2  (    .in(\nand_30.nand_2 ),    .out(\nand_30.and_2 )
  );
  inverter \nand_30.inv_3  (    .in(\nand_30.nand_3 ),    .out(\nand_30.and_3 )
  );
  inverter \nand_30.inv_4  (    .in(\nand_30.nand_4 ),    .out(\nand_30.and_4 )
  );
  nand2 \nand_30.nand2_0  (    .in_0(\in_b<0> ),    .in_1(\in<1> ),    .out(\nand_30.nand_0 )
  );
  nand2 \nand_30.nand2_1  (    .in_0(\nand_30.and_0 ),    .in_1(\in<2> ),    .out(\nand_30.nand_1 )
  );
  nand2 \nand_30.nand2_2  (    .in_0(\nand_30.and_1 ),    .in_1(\in<3> ),    .out(\nand_30.nand_2 )
  );
  nand2 \nand_30.nand2_3  (    .in_0(\nand_30.and_2 ),    .in_1(\in<4> ),    .out(\nand_30.nand_3 )
  );
  nand2 \nand_30.nand2_4  (    .in_0(\nand_30.and_3 ),    .in_1(\in_b<5> ),    .out(\nand_30.nand_4 )
  );
  nand2 \nand_30.nand2_5  (    .in_0(\nand_30.and_4 ),    .in_1(enable),    .out(\nand_30.out )
  );
  inverter \nand_31.inv_0  (    .in(\nand_31.nand_0 ),    .out(\nand_31.and_0 )
  );
  inverter \nand_31.inv_1  (    .in(\nand_31.nand_1 ),    .out(\nand_31.and_1 )
  );
  inverter \nand_31.inv_2  (    .in(\nand_31.nand_2 ),    .out(\nand_31.and_2 )
  );
  inverter \nand_31.inv_3  (    .in(\nand_31.nand_3 ),    .out(\nand_31.and_3 )
  );
  inverter \nand_31.inv_4  (    .in(\nand_31.nand_4 ),    .out(\nand_31.and_4 )
  );
  nand2 \nand_31.nand2_0  (    .in_0(\in<0> ),    .in_1(\in<1> ),    .out(\nand_31.nand_0 )
  );
  nand2 \nand_31.nand2_1  (    .in_0(\nand_31.and_0 ),    .in_1(\in<2> ),    .out(\nand_31.nand_1 )
  );
  nand2 \nand_31.nand2_2  (    .in_0(\nand_31.and_1 ),    .in_1(\in<3> ),    .out(\nand_31.nand_2 )
  );
  nand2 \nand_31.nand2_3  (    .in_0(\nand_31.and_2 ),    .in_1(\in<4> ),    .out(\nand_31.nand_3 )
  );
  nand2 \nand_31.nand2_4  (    .in_0(\nand_31.and_3 ),    .in_1(\in_b<5> ),    .out(\nand_31.nand_4 )
  );
  nand2 \nand_31.nand2_5  (    .in_0(\nand_31.and_4 ),    .in_1(enable),    .out(\nand_31.out )
  );
  inverter \nand_32.inv_0  (    .in(\nand_32.nand_0 ),    .out(\nand_32.and_0 )
  );
  inverter \nand_32.inv_1  (    .in(\nand_32.nand_1 ),    .out(\nand_32.and_1 )
  );
  inverter \nand_32.inv_2  (    .in(\nand_32.nand_2 ),    .out(\nand_32.and_2 )
  );
  inverter \nand_32.inv_3  (    .in(\nand_32.nand_3 ),    .out(\nand_32.and_3 )
  );
  inverter \nand_32.inv_4  (    .in(\nand_32.nand_4 ),    .out(\nand_32.and_4 )
  );
  nand2 \nand_32.nand2_0  (    .in_0(\in_b<0> ),    .in_1(\in_b<1> ),    .out(\nand_32.nand_0 )
  );
  nand2 \nand_32.nand2_1  (    .in_0(\nand_32.and_0 ),    .in_1(\in_b<2> ),    .out(\nand_32.nand_1 )
  );
  nand2 \nand_32.nand2_2  (    .in_0(\nand_32.and_1 ),    .in_1(\in_b<3> ),    .out(\nand_32.nand_2 )
  );
  nand2 \nand_32.nand2_3  (    .in_0(\nand_32.and_2 ),    .in_1(\in_b<4> ),    .out(\nand_32.nand_3 )
  );
  nand2 \nand_32.nand2_4  (    .in_0(\nand_32.and_3 ),    .in_1(\in<5> ),    .out(\nand_32.nand_4 )
  );
  nand2 \nand_32.nand2_5  (    .in_0(\nand_32.and_4 ),    .in_1(enable),    .out(\nand_32.out )
  );
  inverter \nand_33.inv_0  (    .in(\nand_33.nand_0 ),    .out(\nand_33.and_0 )
  );
  inverter \nand_33.inv_1  (    .in(\nand_33.nand_1 ),    .out(\nand_33.and_1 )
  );
  inverter \nand_33.inv_2  (    .in(\nand_33.nand_2 ),    .out(\nand_33.and_2 )
  );
  inverter \nand_33.inv_3  (    .in(\nand_33.nand_3 ),    .out(\nand_33.and_3 )
  );
  inverter \nand_33.inv_4  (    .in(\nand_33.nand_4 ),    .out(\nand_33.and_4 )
  );
  nand2 \nand_33.nand2_0  (    .in_0(\in<0> ),    .in_1(\in_b<1> ),    .out(\nand_33.nand_0 )
  );
  nand2 \nand_33.nand2_1  (    .in_0(\nand_33.and_0 ),    .in_1(\in_b<2> ),    .out(\nand_33.nand_1 )
  );
  nand2 \nand_33.nand2_2  (    .in_0(\nand_33.and_1 ),    .in_1(\in_b<3> ),    .out(\nand_33.nand_2 )
  );
  nand2 \nand_33.nand2_3  (    .in_0(\nand_33.and_2 ),    .in_1(\in_b<4> ),    .out(\nand_33.nand_3 )
  );
  nand2 \nand_33.nand2_4  (    .in_0(\nand_33.and_3 ),    .in_1(\in<5> ),    .out(\nand_33.nand_4 )
  );
  nand2 \nand_33.nand2_5  (    .in_0(\nand_33.and_4 ),    .in_1(enable),    .out(\nand_33.out )
  );
  inverter \nand_34.inv_0  (    .in(\nand_34.nand_0 ),    .out(\nand_34.and_0 )
  );
  inverter \nand_34.inv_1  (    .in(\nand_34.nand_1 ),    .out(\nand_34.and_1 )
  );
  inverter \nand_34.inv_2  (    .in(\nand_34.nand_2 ),    .out(\nand_34.and_2 )
  );
  inverter \nand_34.inv_3  (    .in(\nand_34.nand_3 ),    .out(\nand_34.and_3 )
  );
  inverter \nand_34.inv_4  (    .in(\nand_34.nand_4 ),    .out(\nand_34.and_4 )
  );
  nand2 \nand_34.nand2_0  (    .in_0(\in_b<0> ),    .in_1(\in<1> ),    .out(\nand_34.nand_0 )
  );
  nand2 \nand_34.nand2_1  (    .in_0(\nand_34.and_0 ),    .in_1(\in_b<2> ),    .out(\nand_34.nand_1 )
  );
  nand2 \nand_34.nand2_2  (    .in_0(\nand_34.and_1 ),    .in_1(\in_b<3> ),    .out(\nand_34.nand_2 )
  );
  nand2 \nand_34.nand2_3  (    .in_0(\nand_34.and_2 ),    .in_1(\in_b<4> ),    .out(\nand_34.nand_3 )
  );
  nand2 \nand_34.nand2_4  (    .in_0(\nand_34.and_3 ),    .in_1(\in<5> ),    .out(\nand_34.nand_4 )
  );
  nand2 \nand_34.nand2_5  (    .in_0(\nand_34.and_4 ),    .in_1(enable),    .out(\nand_34.out )
  );
  inverter \nand_35.inv_0  (    .in(\nand_35.nand_0 ),    .out(\nand_35.and_0 )
  );
  inverter \nand_35.inv_1  (    .in(\nand_35.nand_1 ),    .out(\nand_35.and_1 )
  );
  inverter \nand_35.inv_2  (    .in(\nand_35.nand_2 ),    .out(\nand_35.and_2 )
  );
  inverter \nand_35.inv_3  (    .in(\nand_35.nand_3 ),    .out(\nand_35.and_3 )
  );
  inverter \nand_35.inv_4  (    .in(\nand_35.nand_4 ),    .out(\nand_35.and_4 )
  );
  nand2 \nand_35.nand2_0  (    .in_0(\in<0> ),    .in_1(\in<1> ),    .out(\nand_35.nand_0 )
  );
  nand2 \nand_35.nand2_1  (    .in_0(\nand_35.and_0 ),    .in_1(\in_b<2> ),    .out(\nand_35.nand_1 )
  );
  nand2 \nand_35.nand2_2  (    .in_0(\nand_35.and_1 ),    .in_1(\in_b<3> ),    .out(\nand_35.nand_2 )
  );
  nand2 \nand_35.nand2_3  (    .in_0(\nand_35.and_2 ),    .in_1(\in_b<4> ),    .out(\nand_35.nand_3 )
  );
  nand2 \nand_35.nand2_4  (    .in_0(\nand_35.and_3 ),    .in_1(\in<5> ),    .out(\nand_35.nand_4 )
  );
  nand2 \nand_35.nand2_5  (    .in_0(\nand_35.and_4 ),    .in_1(enable),    .out(\nand_35.out )
  );
  inverter \nand_36.inv_0  (    .in(\nand_36.nand_0 ),    .out(\nand_36.and_0 )
  );
  inverter \nand_36.inv_1  (    .in(\nand_36.nand_1 ),    .out(\nand_36.and_1 )
  );
  inverter \nand_36.inv_2  (    .in(\nand_36.nand_2 ),    .out(\nand_36.and_2 )
  );
  inverter \nand_36.inv_3  (    .in(\nand_36.nand_3 ),    .out(\nand_36.and_3 )
  );
  inverter \nand_36.inv_4  (    .in(\nand_36.nand_4 ),    .out(\nand_36.and_4 )
  );
  nand2 \nand_36.nand2_0  (    .in_0(\in_b<0> ),    .in_1(\in_b<1> ),    .out(\nand_36.nand_0 )
  );
  nand2 \nand_36.nand2_1  (    .in_0(\nand_36.and_0 ),    .in_1(\in<2> ),    .out(\nand_36.nand_1 )
  );
  nand2 \nand_36.nand2_2  (    .in_0(\nand_36.and_1 ),    .in_1(\in_b<3> ),    .out(\nand_36.nand_2 )
  );
  nand2 \nand_36.nand2_3  (    .in_0(\nand_36.and_2 ),    .in_1(\in_b<4> ),    .out(\nand_36.nand_3 )
  );
  nand2 \nand_36.nand2_4  (    .in_0(\nand_36.and_3 ),    .in_1(\in<5> ),    .out(\nand_36.nand_4 )
  );
  nand2 \nand_36.nand2_5  (    .in_0(\nand_36.and_4 ),    .in_1(enable),    .out(\nand_36.out )
  );
  inverter \nand_37.inv_0  (    .in(\nand_37.nand_0 ),    .out(\nand_37.and_0 )
  );
  inverter \nand_37.inv_1  (    .in(\nand_37.nand_1 ),    .out(\nand_37.and_1 )
  );
  inverter \nand_37.inv_2  (    .in(\nand_37.nand_2 ),    .out(\nand_37.and_2 )
  );
  inverter \nand_37.inv_3  (    .in(\nand_37.nand_3 ),    .out(\nand_37.and_3 )
  );
  inverter \nand_37.inv_4  (    .in(\nand_37.nand_4 ),    .out(\nand_37.and_4 )
  );
  nand2 \nand_37.nand2_0  (    .in_0(\in<0> ),    .in_1(\in_b<1> ),    .out(\nand_37.nand_0 )
  );
  nand2 \nand_37.nand2_1  (    .in_0(\nand_37.and_0 ),    .in_1(\in<2> ),    .out(\nand_37.nand_1 )
  );
  nand2 \nand_37.nand2_2  (    .in_0(\nand_37.and_1 ),    .in_1(\in_b<3> ),    .out(\nand_37.nand_2 )
  );
  nand2 \nand_37.nand2_3  (    .in_0(\nand_37.and_2 ),    .in_1(\in_b<4> ),    .out(\nand_37.nand_3 )
  );
  nand2 \nand_37.nand2_4  (    .in_0(\nand_37.and_3 ),    .in_1(\in<5> ),    .out(\nand_37.nand_4 )
  );
  nand2 \nand_37.nand2_5  (    .in_0(\nand_37.and_4 ),    .in_1(enable),    .out(\nand_37.out )
  );
  inverter \nand_38.inv_0  (    .in(\nand_38.nand_0 ),    .out(\nand_38.and_0 )
  );
  inverter \nand_38.inv_1  (    .in(\nand_38.nand_1 ),    .out(\nand_38.and_1 )
  );
  inverter \nand_38.inv_2  (    .in(\nand_38.nand_2 ),    .out(\nand_38.and_2 )
  );
  inverter \nand_38.inv_3  (    .in(\nand_38.nand_3 ),    .out(\nand_38.and_3 )
  );
  inverter \nand_38.inv_4  (    .in(\nand_38.nand_4 ),    .out(\nand_38.and_4 )
  );
  nand2 \nand_38.nand2_0  (    .in_0(\in_b<0> ),    .in_1(\in<1> ),    .out(\nand_38.nand_0 )
  );
  nand2 \nand_38.nand2_1  (    .in_0(\nand_38.and_0 ),    .in_1(\in<2> ),    .out(\nand_38.nand_1 )
  );
  nand2 \nand_38.nand2_2  (    .in_0(\nand_38.and_1 ),    .in_1(\in_b<3> ),    .out(\nand_38.nand_2 )
  );
  nand2 \nand_38.nand2_3  (    .in_0(\nand_38.and_2 ),    .in_1(\in_b<4> ),    .out(\nand_38.nand_3 )
  );
  nand2 \nand_38.nand2_4  (    .in_0(\nand_38.and_3 ),    .in_1(\in<5> ),    .out(\nand_38.nand_4 )
  );
  nand2 \nand_38.nand2_5  (    .in_0(\nand_38.and_4 ),    .in_1(enable),    .out(\nand_38.out )
  );
  inverter \nand_39.inv_0  (    .in(\nand_39.nand_0 ),    .out(\nand_39.and_0 )
  );
  inverter \nand_39.inv_1  (    .in(\nand_39.nand_1 ),    .out(\nand_39.and_1 )
  );
  inverter \nand_39.inv_2  (    .in(\nand_39.nand_2 ),    .out(\nand_39.and_2 )
  );
  inverter \nand_39.inv_3  (    .in(\nand_39.nand_3 ),    .out(\nand_39.and_3 )
  );
  inverter \nand_39.inv_4  (    .in(\nand_39.nand_4 ),    .out(\nand_39.and_4 )
  );
  nand2 \nand_39.nand2_0  (    .in_0(\in<0> ),    .in_1(\in<1> ),    .out(\nand_39.nand_0 )
  );
  nand2 \nand_39.nand2_1  (    .in_0(\nand_39.and_0 ),    .in_1(\in<2> ),    .out(\nand_39.nand_1 )
  );
  nand2 \nand_39.nand2_2  (    .in_0(\nand_39.and_1 ),    .in_1(\in_b<3> ),    .out(\nand_39.nand_2 )
  );
  nand2 \nand_39.nand2_3  (    .in_0(\nand_39.and_2 ),    .in_1(\in_b<4> ),    .out(\nand_39.nand_3 )
  );
  nand2 \nand_39.nand2_4  (    .in_0(\nand_39.and_3 ),    .in_1(\in<5> ),    .out(\nand_39.nand_4 )
  );
  nand2 \nand_39.nand2_5  (    .in_0(\nand_39.and_4 ),    .in_1(enable),    .out(\nand_39.out )
  );
  inverter \nand_4.inv_0  (    .in(\nand_4.nand_0 ),    .out(\nand_4.and_0 )
  );
  inverter \nand_4.inv_1  (    .in(\nand_4.nand_1 ),    .out(\nand_4.and_1 )
  );
  inverter \nand_4.inv_2  (    .in(\nand_4.nand_2 ),    .out(\nand_4.and_2 )
  );
  inverter \nand_4.inv_3  (    .in(\nand_4.nand_3 ),    .out(\nand_4.and_3 )
  );
  inverter \nand_4.inv_4  (    .in(\nand_4.nand_4 ),    .out(\nand_4.and_4 )
  );
  nand2 \nand_4.nand2_0  (    .in_0(\in_b<0> ),    .in_1(\in_b<1> ),    .out(\nand_4.nand_0 )
  );
  nand2 \nand_4.nand2_1  (    .in_0(\nand_4.and_0 ),    .in_1(\in<2> ),    .out(\nand_4.nand_1 )
  );
  nand2 \nand_4.nand2_2  (    .in_0(\nand_4.and_1 ),    .in_1(\in_b<3> ),    .out(\nand_4.nand_2 )
  );
  nand2 \nand_4.nand2_3  (    .in_0(\nand_4.and_2 ),    .in_1(\in_b<4> ),    .out(\nand_4.nand_3 )
  );
  nand2 \nand_4.nand2_4  (    .in_0(\nand_4.and_3 ),    .in_1(\in_b<5> ),    .out(\nand_4.nand_4 )
  );
  nand2 \nand_4.nand2_5  (    .in_0(\nand_4.and_4 ),    .in_1(enable),    .out(\nand_4.out )
  );
  inverter \nand_40.inv_0  (    .in(\nand_40.nand_0 ),    .out(\nand_40.and_0 )
  );
  inverter \nand_40.inv_1  (    .in(\nand_40.nand_1 ),    .out(\nand_40.and_1 )
  );
  inverter \nand_40.inv_2  (    .in(\nand_40.nand_2 ),    .out(\nand_40.and_2 )
  );
  inverter \nand_40.inv_3  (    .in(\nand_40.nand_3 ),    .out(\nand_40.and_3 )
  );
  inverter \nand_40.inv_4  (    .in(\nand_40.nand_4 ),    .out(\nand_40.and_4 )
  );
  nand2 \nand_40.nand2_0  (    .in_0(\in_b<0> ),    .in_1(\in_b<1> ),    .out(\nand_40.nand_0 )
  );
  nand2 \nand_40.nand2_1  (    .in_0(\nand_40.and_0 ),    .in_1(\in_b<2> ),    .out(\nand_40.nand_1 )
  );
  nand2 \nand_40.nand2_2  (    .in_0(\nand_40.and_1 ),    .in_1(\in<3> ),    .out(\nand_40.nand_2 )
  );
  nand2 \nand_40.nand2_3  (    .in_0(\nand_40.and_2 ),    .in_1(\in_b<4> ),    .out(\nand_40.nand_3 )
  );
  nand2 \nand_40.nand2_4  (    .in_0(\nand_40.and_3 ),    .in_1(\in<5> ),    .out(\nand_40.nand_4 )
  );
  nand2 \nand_40.nand2_5  (    .in_0(\nand_40.and_4 ),    .in_1(enable),    .out(\nand_40.out )
  );
  inverter \nand_41.inv_0  (    .in(\nand_41.nand_0 ),    .out(\nand_41.and_0 )
  );
  inverter \nand_41.inv_1  (    .in(\nand_41.nand_1 ),    .out(\nand_41.and_1 )
  );
  inverter \nand_41.inv_2  (    .in(\nand_41.nand_2 ),    .out(\nand_41.and_2 )
  );
  inverter \nand_41.inv_3  (    .in(\nand_41.nand_3 ),    .out(\nand_41.and_3 )
  );
  inverter \nand_41.inv_4  (    .in(\nand_41.nand_4 ),    .out(\nand_41.and_4 )
  );
  nand2 \nand_41.nand2_0  (    .in_0(\in<0> ),    .in_1(\in_b<1> ),    .out(\nand_41.nand_0 )
  );
  nand2 \nand_41.nand2_1  (    .in_0(\nand_41.and_0 ),    .in_1(\in_b<2> ),    .out(\nand_41.nand_1 )
  );
  nand2 \nand_41.nand2_2  (    .in_0(\nand_41.and_1 ),    .in_1(\in<3> ),    .out(\nand_41.nand_2 )
  );
  nand2 \nand_41.nand2_3  (    .in_0(\nand_41.and_2 ),    .in_1(\in_b<4> ),    .out(\nand_41.nand_3 )
  );
  nand2 \nand_41.nand2_4  (    .in_0(\nand_41.and_3 ),    .in_1(\in<5> ),    .out(\nand_41.nand_4 )
  );
  nand2 \nand_41.nand2_5  (    .in_0(\nand_41.and_4 ),    .in_1(enable),    .out(\nand_41.out )
  );
  inverter \nand_42.inv_0  (    .in(\nand_42.nand_0 ),    .out(\nand_42.and_0 )
  );
  inverter \nand_42.inv_1  (    .in(\nand_42.nand_1 ),    .out(\nand_42.and_1 )
  );
  inverter \nand_42.inv_2  (    .in(\nand_42.nand_2 ),    .out(\nand_42.and_2 )
  );
  inverter \nand_42.inv_3  (    .in(\nand_42.nand_3 ),    .out(\nand_42.and_3 )
  );
  inverter \nand_42.inv_4  (    .in(\nand_42.nand_4 ),    .out(\nand_42.and_4 )
  );
  nand2 \nand_42.nand2_0  (    .in_0(\in_b<0> ),    .in_1(\in<1> ),    .out(\nand_42.nand_0 )
  );
  nand2 \nand_42.nand2_1  (    .in_0(\nand_42.and_0 ),    .in_1(\in_b<2> ),    .out(\nand_42.nand_1 )
  );
  nand2 \nand_42.nand2_2  (    .in_0(\nand_42.and_1 ),    .in_1(\in<3> ),    .out(\nand_42.nand_2 )
  );
  nand2 \nand_42.nand2_3  (    .in_0(\nand_42.and_2 ),    .in_1(\in_b<4> ),    .out(\nand_42.nand_3 )
  );
  nand2 \nand_42.nand2_4  (    .in_0(\nand_42.and_3 ),    .in_1(\in<5> ),    .out(\nand_42.nand_4 )
  );
  nand2 \nand_42.nand2_5  (    .in_0(\nand_42.and_4 ),    .in_1(enable),    .out(\nand_42.out )
  );
  inverter \nand_43.inv_0  (    .in(\nand_43.nand_0 ),    .out(\nand_43.and_0 )
  );
  inverter \nand_43.inv_1  (    .in(\nand_43.nand_1 ),    .out(\nand_43.and_1 )
  );
  inverter \nand_43.inv_2  (    .in(\nand_43.nand_2 ),    .out(\nand_43.and_2 )
  );
  inverter \nand_43.inv_3  (    .in(\nand_43.nand_3 ),    .out(\nand_43.and_3 )
  );
  inverter \nand_43.inv_4  (    .in(\nand_43.nand_4 ),    .out(\nand_43.and_4 )
  );
  nand2 \nand_43.nand2_0  (    .in_0(\in<0> ),    .in_1(\in<1> ),    .out(\nand_43.nand_0 )
  );
  nand2 \nand_43.nand2_1  (    .in_0(\nand_43.and_0 ),    .in_1(\in_b<2> ),    .out(\nand_43.nand_1 )
  );
  nand2 \nand_43.nand2_2  (    .in_0(\nand_43.and_1 ),    .in_1(\in<3> ),    .out(\nand_43.nand_2 )
  );
  nand2 \nand_43.nand2_3  (    .in_0(\nand_43.and_2 ),    .in_1(\in_b<4> ),    .out(\nand_43.nand_3 )
  );
  nand2 \nand_43.nand2_4  (    .in_0(\nand_43.and_3 ),    .in_1(\in<5> ),    .out(\nand_43.nand_4 )
  );
  nand2 \nand_43.nand2_5  (    .in_0(\nand_43.and_4 ),    .in_1(enable),    .out(\nand_43.out )
  );
  inverter \nand_44.inv_0  (    .in(\nand_44.nand_0 ),    .out(\nand_44.and_0 )
  );
  inverter \nand_44.inv_1  (    .in(\nand_44.nand_1 ),    .out(\nand_44.and_1 )
  );
  inverter \nand_44.inv_2  (    .in(\nand_44.nand_2 ),    .out(\nand_44.and_2 )
  );
  inverter \nand_44.inv_3  (    .in(\nand_44.nand_3 ),    .out(\nand_44.and_3 )
  );
  inverter \nand_44.inv_4  (    .in(\nand_44.nand_4 ),    .out(\nand_44.and_4 )
  );
  nand2 \nand_44.nand2_0  (    .in_0(\in_b<0> ),    .in_1(\in_b<1> ),    .out(\nand_44.nand_0 )
  );
  nand2 \nand_44.nand2_1  (    .in_0(\nand_44.and_0 ),    .in_1(\in<2> ),    .out(\nand_44.nand_1 )
  );
  nand2 \nand_44.nand2_2  (    .in_0(\nand_44.and_1 ),    .in_1(\in<3> ),    .out(\nand_44.nand_2 )
  );
  nand2 \nand_44.nand2_3  (    .in_0(\nand_44.and_2 ),    .in_1(\in_b<4> ),    .out(\nand_44.nand_3 )
  );
  nand2 \nand_44.nand2_4  (    .in_0(\nand_44.and_3 ),    .in_1(\in<5> ),    .out(\nand_44.nand_4 )
  );
  nand2 \nand_44.nand2_5  (    .in_0(\nand_44.and_4 ),    .in_1(enable),    .out(\nand_44.out )
  );
  inverter \nand_45.inv_0  (    .in(\nand_45.nand_0 ),    .out(\nand_45.and_0 )
  );
  inverter \nand_45.inv_1  (    .in(\nand_45.nand_1 ),    .out(\nand_45.and_1 )
  );
  inverter \nand_45.inv_2  (    .in(\nand_45.nand_2 ),    .out(\nand_45.and_2 )
  );
  inverter \nand_45.inv_3  (    .in(\nand_45.nand_3 ),    .out(\nand_45.and_3 )
  );
  inverter \nand_45.inv_4  (    .in(\nand_45.nand_4 ),    .out(\nand_45.and_4 )
  );
  nand2 \nand_45.nand2_0  (    .in_0(\in<0> ),    .in_1(\in_b<1> ),    .out(\nand_45.nand_0 )
  );
  nand2 \nand_45.nand2_1  (    .in_0(\nand_45.and_0 ),    .in_1(\in<2> ),    .out(\nand_45.nand_1 )
  );
  nand2 \nand_45.nand2_2  (    .in_0(\nand_45.and_1 ),    .in_1(\in<3> ),    .out(\nand_45.nand_2 )
  );
  nand2 \nand_45.nand2_3  (    .in_0(\nand_45.and_2 ),    .in_1(\in_b<4> ),    .out(\nand_45.nand_3 )
  );
  nand2 \nand_45.nand2_4  (    .in_0(\nand_45.and_3 ),    .in_1(\in<5> ),    .out(\nand_45.nand_4 )
  );
  nand2 \nand_45.nand2_5  (    .in_0(\nand_45.and_4 ),    .in_1(enable),    .out(\nand_45.out )
  );
  inverter \nand_46.inv_0  (    .in(\nand_46.nand_0 ),    .out(\nand_46.and_0 )
  );
  inverter \nand_46.inv_1  (    .in(\nand_46.nand_1 ),    .out(\nand_46.and_1 )
  );
  inverter \nand_46.inv_2  (    .in(\nand_46.nand_2 ),    .out(\nand_46.and_2 )
  );
  inverter \nand_46.inv_3  (    .in(\nand_46.nand_3 ),    .out(\nand_46.and_3 )
  );
  inverter \nand_46.inv_4  (    .in(\nand_46.nand_4 ),    .out(\nand_46.and_4 )
  );
  nand2 \nand_46.nand2_0  (    .in_0(\in_b<0> ),    .in_1(\in<1> ),    .out(\nand_46.nand_0 )
  );
  nand2 \nand_46.nand2_1  (    .in_0(\nand_46.and_0 ),    .in_1(\in<2> ),    .out(\nand_46.nand_1 )
  );
  nand2 \nand_46.nand2_2  (    .in_0(\nand_46.and_1 ),    .in_1(\in<3> ),    .out(\nand_46.nand_2 )
  );
  nand2 \nand_46.nand2_3  (    .in_0(\nand_46.and_2 ),    .in_1(\in_b<4> ),    .out(\nand_46.nand_3 )
  );
  nand2 \nand_46.nand2_4  (    .in_0(\nand_46.and_3 ),    .in_1(\in<5> ),    .out(\nand_46.nand_4 )
  );
  nand2 \nand_46.nand2_5  (    .in_0(\nand_46.and_4 ),    .in_1(enable),    .out(\nand_46.out )
  );
  inverter \nand_47.inv_0  (    .in(\nand_47.nand_0 ),    .out(\nand_47.and_0 )
  );
  inverter \nand_47.inv_1  (    .in(\nand_47.nand_1 ),    .out(\nand_47.and_1 )
  );
  inverter \nand_47.inv_2  (    .in(\nand_47.nand_2 ),    .out(\nand_47.and_2 )
  );
  inverter \nand_47.inv_3  (    .in(\nand_47.nand_3 ),    .out(\nand_47.and_3 )
  );
  inverter \nand_47.inv_4  (    .in(\nand_47.nand_4 ),    .out(\nand_47.and_4 )
  );
  nand2 \nand_47.nand2_0  (    .in_0(\in<0> ),    .in_1(\in<1> ),    .out(\nand_47.nand_0 )
  );
  nand2 \nand_47.nand2_1  (    .in_0(\nand_47.and_0 ),    .in_1(\in<2> ),    .out(\nand_47.nand_1 )
  );
  nand2 \nand_47.nand2_2  (    .in_0(\nand_47.and_1 ),    .in_1(\in<3> ),    .out(\nand_47.nand_2 )
  );
  nand2 \nand_47.nand2_3  (    .in_0(\nand_47.and_2 ),    .in_1(\in_b<4> ),    .out(\nand_47.nand_3 )
  );
  nand2 \nand_47.nand2_4  (    .in_0(\nand_47.and_3 ),    .in_1(\in<5> ),    .out(\nand_47.nand_4 )
  );
  nand2 \nand_47.nand2_5  (    .in_0(\nand_47.and_4 ),    .in_1(enable),    .out(\nand_47.out )
  );
  inverter \nand_48.inv_0  (    .in(\nand_48.nand_0 ),    .out(\nand_48.and_0 )
  );
  inverter \nand_48.inv_1  (    .in(\nand_48.nand_1 ),    .out(\nand_48.and_1 )
  );
  inverter \nand_48.inv_2  (    .in(\nand_48.nand_2 ),    .out(\nand_48.and_2 )
  );
  inverter \nand_48.inv_3  (    .in(\nand_48.nand_3 ),    .out(\nand_48.and_3 )
  );
  inverter \nand_48.inv_4  (    .in(\nand_48.nand_4 ),    .out(\nand_48.and_4 )
  );
  nand2 \nand_48.nand2_0  (    .in_0(\in_b<0> ),    .in_1(\in_b<1> ),    .out(\nand_48.nand_0 )
  );
  nand2 \nand_48.nand2_1  (    .in_0(\nand_48.and_0 ),    .in_1(\in_b<2> ),    .out(\nand_48.nand_1 )
  );
  nand2 \nand_48.nand2_2  (    .in_0(\nand_48.and_1 ),    .in_1(\in_b<3> ),    .out(\nand_48.nand_2 )
  );
  nand2 \nand_48.nand2_3  (    .in_0(\nand_48.and_2 ),    .in_1(\in<4> ),    .out(\nand_48.nand_3 )
  );
  nand2 \nand_48.nand2_4  (    .in_0(\nand_48.and_3 ),    .in_1(\in<5> ),    .out(\nand_48.nand_4 )
  );
  nand2 \nand_48.nand2_5  (    .in_0(\nand_48.and_4 ),    .in_1(enable),    .out(\nand_48.out )
  );
  inverter \nand_49.inv_0  (    .in(\nand_49.nand_0 ),    .out(\nand_49.and_0 )
  );
  inverter \nand_49.inv_1  (    .in(\nand_49.nand_1 ),    .out(\nand_49.and_1 )
  );
  inverter \nand_49.inv_2  (    .in(\nand_49.nand_2 ),    .out(\nand_49.and_2 )
  );
  inverter \nand_49.inv_3  (    .in(\nand_49.nand_3 ),    .out(\nand_49.and_3 )
  );
  inverter \nand_49.inv_4  (    .in(\nand_49.nand_4 ),    .out(\nand_49.and_4 )
  );
  nand2 \nand_49.nand2_0  (    .in_0(\in<0> ),    .in_1(\in_b<1> ),    .out(\nand_49.nand_0 )
  );
  nand2 \nand_49.nand2_1  (    .in_0(\nand_49.and_0 ),    .in_1(\in_b<2> ),    .out(\nand_49.nand_1 )
  );
  nand2 \nand_49.nand2_2  (    .in_0(\nand_49.and_1 ),    .in_1(\in_b<3> ),    .out(\nand_49.nand_2 )
  );
  nand2 \nand_49.nand2_3  (    .in_0(\nand_49.and_2 ),    .in_1(\in<4> ),    .out(\nand_49.nand_3 )
  );
  nand2 \nand_49.nand2_4  (    .in_0(\nand_49.and_3 ),    .in_1(\in<5> ),    .out(\nand_49.nand_4 )
  );
  nand2 \nand_49.nand2_5  (    .in_0(\nand_49.and_4 ),    .in_1(enable),    .out(\nand_49.out )
  );
  inverter \nand_5.inv_0  (    .in(\nand_5.nand_0 ),    .out(\nand_5.and_0 )
  );
  inverter \nand_5.inv_1  (    .in(\nand_5.nand_1 ),    .out(\nand_5.and_1 )
  );
  inverter \nand_5.inv_2  (    .in(\nand_5.nand_2 ),    .out(\nand_5.and_2 )
  );
  inverter \nand_5.inv_3  (    .in(\nand_5.nand_3 ),    .out(\nand_5.and_3 )
  );
  inverter \nand_5.inv_4  (    .in(\nand_5.nand_4 ),    .out(\nand_5.and_4 )
  );
  nand2 \nand_5.nand2_0  (    .in_0(\in<0> ),    .in_1(\in_b<1> ),    .out(\nand_5.nand_0 )
  );
  nand2 \nand_5.nand2_1  (    .in_0(\nand_5.and_0 ),    .in_1(\in<2> ),    .out(\nand_5.nand_1 )
  );
  nand2 \nand_5.nand2_2  (    .in_0(\nand_5.and_1 ),    .in_1(\in_b<3> ),    .out(\nand_5.nand_2 )
  );
  nand2 \nand_5.nand2_3  (    .in_0(\nand_5.and_2 ),    .in_1(\in_b<4> ),    .out(\nand_5.nand_3 )
  );
  nand2 \nand_5.nand2_4  (    .in_0(\nand_5.and_3 ),    .in_1(\in_b<5> ),    .out(\nand_5.nand_4 )
  );
  nand2 \nand_5.nand2_5  (    .in_0(\nand_5.and_4 ),    .in_1(enable),    .out(\nand_5.out )
  );
  inverter \nand_50.inv_0  (    .in(\nand_50.nand_0 ),    .out(\nand_50.and_0 )
  );
  inverter \nand_50.inv_1  (    .in(\nand_50.nand_1 ),    .out(\nand_50.and_1 )
  );
  inverter \nand_50.inv_2  (    .in(\nand_50.nand_2 ),    .out(\nand_50.and_2 )
  );
  inverter \nand_50.inv_3  (    .in(\nand_50.nand_3 ),    .out(\nand_50.and_3 )
  );
  inverter \nand_50.inv_4  (    .in(\nand_50.nand_4 ),    .out(\nand_50.and_4 )
  );
  nand2 \nand_50.nand2_0  (    .in_0(\in_b<0> ),    .in_1(\in<1> ),    .out(\nand_50.nand_0 )
  );
  nand2 \nand_50.nand2_1  (    .in_0(\nand_50.and_0 ),    .in_1(\in_b<2> ),    .out(\nand_50.nand_1 )
  );
  nand2 \nand_50.nand2_2  (    .in_0(\nand_50.and_1 ),    .in_1(\in_b<3> ),    .out(\nand_50.nand_2 )
  );
  nand2 \nand_50.nand2_3  (    .in_0(\nand_50.and_2 ),    .in_1(\in<4> ),    .out(\nand_50.nand_3 )
  );
  nand2 \nand_50.nand2_4  (    .in_0(\nand_50.and_3 ),    .in_1(\in<5> ),    .out(\nand_50.nand_4 )
  );
  nand2 \nand_50.nand2_5  (    .in_0(\nand_50.and_4 ),    .in_1(enable),    .out(\nand_50.out )
  );
  inverter \nand_51.inv_0  (    .in(\nand_51.nand_0 ),    .out(\nand_51.and_0 )
  );
  inverter \nand_51.inv_1  (    .in(\nand_51.nand_1 ),    .out(\nand_51.and_1 )
  );
  inverter \nand_51.inv_2  (    .in(\nand_51.nand_2 ),    .out(\nand_51.and_2 )
  );
  inverter \nand_51.inv_3  (    .in(\nand_51.nand_3 ),    .out(\nand_51.and_3 )
  );
  inverter \nand_51.inv_4  (    .in(\nand_51.nand_4 ),    .out(\nand_51.and_4 )
  );
  nand2 \nand_51.nand2_0  (    .in_0(\in<0> ),    .in_1(\in<1> ),    .out(\nand_51.nand_0 )
  );
  nand2 \nand_51.nand2_1  (    .in_0(\nand_51.and_0 ),    .in_1(\in_b<2> ),    .out(\nand_51.nand_1 )
  );
  nand2 \nand_51.nand2_2  (    .in_0(\nand_51.and_1 ),    .in_1(\in_b<3> ),    .out(\nand_51.nand_2 )
  );
  nand2 \nand_51.nand2_3  (    .in_0(\nand_51.and_2 ),    .in_1(\in<4> ),    .out(\nand_51.nand_3 )
  );
  nand2 \nand_51.nand2_4  (    .in_0(\nand_51.and_3 ),    .in_1(\in<5> ),    .out(\nand_51.nand_4 )
  );
  nand2 \nand_51.nand2_5  (    .in_0(\nand_51.and_4 ),    .in_1(enable),    .out(\nand_51.out )
  );
  inverter \nand_52.inv_0  (    .in(\nand_52.nand_0 ),    .out(\nand_52.and_0 )
  );
  inverter \nand_52.inv_1  (    .in(\nand_52.nand_1 ),    .out(\nand_52.and_1 )
  );
  inverter \nand_52.inv_2  (    .in(\nand_52.nand_2 ),    .out(\nand_52.and_2 )
  );
  inverter \nand_52.inv_3  (    .in(\nand_52.nand_3 ),    .out(\nand_52.and_3 )
  );
  inverter \nand_52.inv_4  (    .in(\nand_52.nand_4 ),    .out(\nand_52.and_4 )
  );
  nand2 \nand_52.nand2_0  (    .in_0(\in_b<0> ),    .in_1(\in_b<1> ),    .out(\nand_52.nand_0 )
  );
  nand2 \nand_52.nand2_1  (    .in_0(\nand_52.and_0 ),    .in_1(\in<2> ),    .out(\nand_52.nand_1 )
  );
  nand2 \nand_52.nand2_2  (    .in_0(\nand_52.and_1 ),    .in_1(\in_b<3> ),    .out(\nand_52.nand_2 )
  );
  nand2 \nand_52.nand2_3  (    .in_0(\nand_52.and_2 ),    .in_1(\in<4> ),    .out(\nand_52.nand_3 )
  );
  nand2 \nand_52.nand2_4  (    .in_0(\nand_52.and_3 ),    .in_1(\in<5> ),    .out(\nand_52.nand_4 )
  );
  nand2 \nand_52.nand2_5  (    .in_0(\nand_52.and_4 ),    .in_1(enable),    .out(\nand_52.out )
  );
  inverter \nand_53.inv_0  (    .in(\nand_53.nand_0 ),    .out(\nand_53.and_0 )
  );
  inverter \nand_53.inv_1  (    .in(\nand_53.nand_1 ),    .out(\nand_53.and_1 )
  );
  inverter \nand_53.inv_2  (    .in(\nand_53.nand_2 ),    .out(\nand_53.and_2 )
  );
  inverter \nand_53.inv_3  (    .in(\nand_53.nand_3 ),    .out(\nand_53.and_3 )
  );
  inverter \nand_53.inv_4  (    .in(\nand_53.nand_4 ),    .out(\nand_53.and_4 )
  );
  nand2 \nand_53.nand2_0  (    .in_0(\in<0> ),    .in_1(\in_b<1> ),    .out(\nand_53.nand_0 )
  );
  nand2 \nand_53.nand2_1  (    .in_0(\nand_53.and_0 ),    .in_1(\in<2> ),    .out(\nand_53.nand_1 )
  );
  nand2 \nand_53.nand2_2  (    .in_0(\nand_53.and_1 ),    .in_1(\in_b<3> ),    .out(\nand_53.nand_2 )
  );
  nand2 \nand_53.nand2_3  (    .in_0(\nand_53.and_2 ),    .in_1(\in<4> ),    .out(\nand_53.nand_3 )
  );
  nand2 \nand_53.nand2_4  (    .in_0(\nand_53.and_3 ),    .in_1(\in<5> ),    .out(\nand_53.nand_4 )
  );
  nand2 \nand_53.nand2_5  (    .in_0(\nand_53.and_4 ),    .in_1(enable),    .out(\nand_53.out )
  );
  inverter \nand_54.inv_0  (    .in(\nand_54.nand_0 ),    .out(\nand_54.and_0 )
  );
  inverter \nand_54.inv_1  (    .in(\nand_54.nand_1 ),    .out(\nand_54.and_1 )
  );
  inverter \nand_54.inv_2  (    .in(\nand_54.nand_2 ),    .out(\nand_54.and_2 )
  );
  inverter \nand_54.inv_3  (    .in(\nand_54.nand_3 ),    .out(\nand_54.and_3 )
  );
  inverter \nand_54.inv_4  (    .in(\nand_54.nand_4 ),    .out(\nand_54.and_4 )
  );
  nand2 \nand_54.nand2_0  (    .in_0(\in_b<0> ),    .in_1(\in<1> ),    .out(\nand_54.nand_0 )
  );
  nand2 \nand_54.nand2_1  (    .in_0(\nand_54.and_0 ),    .in_1(\in<2> ),    .out(\nand_54.nand_1 )
  );
  nand2 \nand_54.nand2_2  (    .in_0(\nand_54.and_1 ),    .in_1(\in_b<3> ),    .out(\nand_54.nand_2 )
  );
  nand2 \nand_54.nand2_3  (    .in_0(\nand_54.and_2 ),    .in_1(\in<4> ),    .out(\nand_54.nand_3 )
  );
  nand2 \nand_54.nand2_4  (    .in_0(\nand_54.and_3 ),    .in_1(\in<5> ),    .out(\nand_54.nand_4 )
  );
  nand2 \nand_54.nand2_5  (    .in_0(\nand_54.and_4 ),    .in_1(enable),    .out(\nand_54.out )
  );
  inverter \nand_55.inv_0  (    .in(\nand_55.nand_0 ),    .out(\nand_55.and_0 )
  );
  inverter \nand_55.inv_1  (    .in(\nand_55.nand_1 ),    .out(\nand_55.and_1 )
  );
  inverter \nand_55.inv_2  (    .in(\nand_55.nand_2 ),    .out(\nand_55.and_2 )
  );
  inverter \nand_55.inv_3  (    .in(\nand_55.nand_3 ),    .out(\nand_55.and_3 )
  );
  inverter \nand_55.inv_4  (    .in(\nand_55.nand_4 ),    .out(\nand_55.and_4 )
  );
  nand2 \nand_55.nand2_0  (    .in_0(\in<0> ),    .in_1(\in<1> ),    .out(\nand_55.nand_0 )
  );
  nand2 \nand_55.nand2_1  (    .in_0(\nand_55.and_0 ),    .in_1(\in<2> ),    .out(\nand_55.nand_1 )
  );
  nand2 \nand_55.nand2_2  (    .in_0(\nand_55.and_1 ),    .in_1(\in_b<3> ),    .out(\nand_55.nand_2 )
  );
  nand2 \nand_55.nand2_3  (    .in_0(\nand_55.and_2 ),    .in_1(\in<4> ),    .out(\nand_55.nand_3 )
  );
  nand2 \nand_55.nand2_4  (    .in_0(\nand_55.and_3 ),    .in_1(\in<5> ),    .out(\nand_55.nand_4 )
  );
  nand2 \nand_55.nand2_5  (    .in_0(\nand_55.and_4 ),    .in_1(enable),    .out(\nand_55.out )
  );
  inverter \nand_56.inv_0  (    .in(\nand_56.nand_0 ),    .out(\nand_56.and_0 )
  );
  inverter \nand_56.inv_1  (    .in(\nand_56.nand_1 ),    .out(\nand_56.and_1 )
  );
  inverter \nand_56.inv_2  (    .in(\nand_56.nand_2 ),    .out(\nand_56.and_2 )
  );
  inverter \nand_56.inv_3  (    .in(\nand_56.nand_3 ),    .out(\nand_56.and_3 )
  );
  inverter \nand_56.inv_4  (    .in(\nand_56.nand_4 ),    .out(\nand_56.and_4 )
  );
  nand2 \nand_56.nand2_0  (    .in_0(\in_b<0> ),    .in_1(\in_b<1> ),    .out(\nand_56.nand_0 )
  );
  nand2 \nand_56.nand2_1  (    .in_0(\nand_56.and_0 ),    .in_1(\in_b<2> ),    .out(\nand_56.nand_1 )
  );
  nand2 \nand_56.nand2_2  (    .in_0(\nand_56.and_1 ),    .in_1(\in<3> ),    .out(\nand_56.nand_2 )
  );
  nand2 \nand_56.nand2_3  (    .in_0(\nand_56.and_2 ),    .in_1(\in<4> ),    .out(\nand_56.nand_3 )
  );
  nand2 \nand_56.nand2_4  (    .in_0(\nand_56.and_3 ),    .in_1(\in<5> ),    .out(\nand_56.nand_4 )
  );
  nand2 \nand_56.nand2_5  (    .in_0(\nand_56.and_4 ),    .in_1(enable),    .out(\nand_56.out )
  );
  inverter \nand_57.inv_0  (    .in(\nand_57.nand_0 ),    .out(\nand_57.and_0 )
  );
  inverter \nand_57.inv_1  (    .in(\nand_57.nand_1 ),    .out(\nand_57.and_1 )
  );
  inverter \nand_57.inv_2  (    .in(\nand_57.nand_2 ),    .out(\nand_57.and_2 )
  );
  inverter \nand_57.inv_3  (    .in(\nand_57.nand_3 ),    .out(\nand_57.and_3 )
  );
  inverter \nand_57.inv_4  (    .in(\nand_57.nand_4 ),    .out(\nand_57.and_4 )
  );
  nand2 \nand_57.nand2_0  (    .in_0(\in<0> ),    .in_1(\in_b<1> ),    .out(\nand_57.nand_0 )
  );
  nand2 \nand_57.nand2_1  (    .in_0(\nand_57.and_0 ),    .in_1(\in_b<2> ),    .out(\nand_57.nand_1 )
  );
  nand2 \nand_57.nand2_2  (    .in_0(\nand_57.and_1 ),    .in_1(\in<3> ),    .out(\nand_57.nand_2 )
  );
  nand2 \nand_57.nand2_3  (    .in_0(\nand_57.and_2 ),    .in_1(\in<4> ),    .out(\nand_57.nand_3 )
  );
  nand2 \nand_57.nand2_4  (    .in_0(\nand_57.and_3 ),    .in_1(\in<5> ),    .out(\nand_57.nand_4 )
  );
  nand2 \nand_57.nand2_5  (    .in_0(\nand_57.and_4 ),    .in_1(enable),    .out(\nand_57.out )
  );
  inverter \nand_58.inv_0  (    .in(\nand_58.nand_0 ),    .out(\nand_58.and_0 )
  );
  inverter \nand_58.inv_1  (    .in(\nand_58.nand_1 ),    .out(\nand_58.and_1 )
  );
  inverter \nand_58.inv_2  (    .in(\nand_58.nand_2 ),    .out(\nand_58.and_2 )
  );
  inverter \nand_58.inv_3  (    .in(\nand_58.nand_3 ),    .out(\nand_58.and_3 )
  );
  inverter \nand_58.inv_4  (    .in(\nand_58.nand_4 ),    .out(\nand_58.and_4 )
  );
  nand2 \nand_58.nand2_0  (    .in_0(\in_b<0> ),    .in_1(\in<1> ),    .out(\nand_58.nand_0 )
  );
  nand2 \nand_58.nand2_1  (    .in_0(\nand_58.and_0 ),    .in_1(\in_b<2> ),    .out(\nand_58.nand_1 )
  );
  nand2 \nand_58.nand2_2  (    .in_0(\nand_58.and_1 ),    .in_1(\in<3> ),    .out(\nand_58.nand_2 )
  );
  nand2 \nand_58.nand2_3  (    .in_0(\nand_58.and_2 ),    .in_1(\in<4> ),    .out(\nand_58.nand_3 )
  );
  nand2 \nand_58.nand2_4  (    .in_0(\nand_58.and_3 ),    .in_1(\in<5> ),    .out(\nand_58.nand_4 )
  );
  nand2 \nand_58.nand2_5  (    .in_0(\nand_58.and_4 ),    .in_1(enable),    .out(\nand_58.out )
  );
  inverter \nand_59.inv_0  (    .in(\nand_59.nand_0 ),    .out(\nand_59.and_0 )
  );
  inverter \nand_59.inv_1  (    .in(\nand_59.nand_1 ),    .out(\nand_59.and_1 )
  );
  inverter \nand_59.inv_2  (    .in(\nand_59.nand_2 ),    .out(\nand_59.and_2 )
  );
  inverter \nand_59.inv_3  (    .in(\nand_59.nand_3 ),    .out(\nand_59.and_3 )
  );
  inverter \nand_59.inv_4  (    .in(\nand_59.nand_4 ),    .out(\nand_59.and_4 )
  );
  nand2 \nand_59.nand2_0  (    .in_0(\in<0> ),    .in_1(\in<1> ),    .out(\nand_59.nand_0 )
  );
  nand2 \nand_59.nand2_1  (    .in_0(\nand_59.and_0 ),    .in_1(\in_b<2> ),    .out(\nand_59.nand_1 )
  );
  nand2 \nand_59.nand2_2  (    .in_0(\nand_59.and_1 ),    .in_1(\in<3> ),    .out(\nand_59.nand_2 )
  );
  nand2 \nand_59.nand2_3  (    .in_0(\nand_59.and_2 ),    .in_1(\in<4> ),    .out(\nand_59.nand_3 )
  );
  nand2 \nand_59.nand2_4  (    .in_0(\nand_59.and_3 ),    .in_1(\in<5> ),    .out(\nand_59.nand_4 )
  );
  nand2 \nand_59.nand2_5  (    .in_0(\nand_59.and_4 ),    .in_1(enable),    .out(\nand_59.out )
  );
  inverter \nand_6.inv_0  (    .in(\nand_6.nand_0 ),    .out(\nand_6.and_0 )
  );
  inverter \nand_6.inv_1  (    .in(\nand_6.nand_1 ),    .out(\nand_6.and_1 )
  );
  inverter \nand_6.inv_2  (    .in(\nand_6.nand_2 ),    .out(\nand_6.and_2 )
  );
  inverter \nand_6.inv_3  (    .in(\nand_6.nand_3 ),    .out(\nand_6.and_3 )
  );
  inverter \nand_6.inv_4  (    .in(\nand_6.nand_4 ),    .out(\nand_6.and_4 )
  );
  nand2 \nand_6.nand2_0  (    .in_0(\in_b<0> ),    .in_1(\in<1> ),    .out(\nand_6.nand_0 )
  );
  nand2 \nand_6.nand2_1  (    .in_0(\nand_6.and_0 ),    .in_1(\in<2> ),    .out(\nand_6.nand_1 )
  );
  nand2 \nand_6.nand2_2  (    .in_0(\nand_6.and_1 ),    .in_1(\in_b<3> ),    .out(\nand_6.nand_2 )
  );
  nand2 \nand_6.nand2_3  (    .in_0(\nand_6.and_2 ),    .in_1(\in_b<4> ),    .out(\nand_6.nand_3 )
  );
  nand2 \nand_6.nand2_4  (    .in_0(\nand_6.and_3 ),    .in_1(\in_b<5> ),    .out(\nand_6.nand_4 )
  );
  nand2 \nand_6.nand2_5  (    .in_0(\nand_6.and_4 ),    .in_1(enable),    .out(\nand_6.out )
  );
  inverter \nand_60.inv_0  (    .in(\nand_60.nand_0 ),    .out(\nand_60.and_0 )
  );
  inverter \nand_60.inv_1  (    .in(\nand_60.nand_1 ),    .out(\nand_60.and_1 )
  );
  inverter \nand_60.inv_2  (    .in(\nand_60.nand_2 ),    .out(\nand_60.and_2 )
  );
  inverter \nand_60.inv_3  (    .in(\nand_60.nand_3 ),    .out(\nand_60.and_3 )
  );
  inverter \nand_60.inv_4  (    .in(\nand_60.nand_4 ),    .out(\nand_60.and_4 )
  );
  nand2 \nand_60.nand2_0  (    .in_0(\in_b<0> ),    .in_1(\in_b<1> ),    .out(\nand_60.nand_0 )
  );
  nand2 \nand_60.nand2_1  (    .in_0(\nand_60.and_0 ),    .in_1(\in<2> ),    .out(\nand_60.nand_1 )
  );
  nand2 \nand_60.nand2_2  (    .in_0(\nand_60.and_1 ),    .in_1(\in<3> ),    .out(\nand_60.nand_2 )
  );
  nand2 \nand_60.nand2_3  (    .in_0(\nand_60.and_2 ),    .in_1(\in<4> ),    .out(\nand_60.nand_3 )
  );
  nand2 \nand_60.nand2_4  (    .in_0(\nand_60.and_3 ),    .in_1(\in<5> ),    .out(\nand_60.nand_4 )
  );
  nand2 \nand_60.nand2_5  (    .in_0(\nand_60.and_4 ),    .in_1(enable),    .out(\nand_60.out )
  );
  inverter \nand_61.inv_0  (    .in(\nand_61.nand_0 ),    .out(\nand_61.and_0 )
  );
  inverter \nand_61.inv_1  (    .in(\nand_61.nand_1 ),    .out(\nand_61.and_1 )
  );
  inverter \nand_61.inv_2  (    .in(\nand_61.nand_2 ),    .out(\nand_61.and_2 )
  );
  inverter \nand_61.inv_3  (    .in(\nand_61.nand_3 ),    .out(\nand_61.and_3 )
  );
  inverter \nand_61.inv_4  (    .in(\nand_61.nand_4 ),    .out(\nand_61.and_4 )
  );
  nand2 \nand_61.nand2_0  (    .in_0(\in<0> ),    .in_1(\in_b<1> ),    .out(\nand_61.nand_0 )
  );
  nand2 \nand_61.nand2_1  (    .in_0(\nand_61.and_0 ),    .in_1(\in<2> ),    .out(\nand_61.nand_1 )
  );
  nand2 \nand_61.nand2_2  (    .in_0(\nand_61.and_1 ),    .in_1(\in<3> ),    .out(\nand_61.nand_2 )
  );
  nand2 \nand_61.nand2_3  (    .in_0(\nand_61.and_2 ),    .in_1(\in<4> ),    .out(\nand_61.nand_3 )
  );
  nand2 \nand_61.nand2_4  (    .in_0(\nand_61.and_3 ),    .in_1(\in<5> ),    .out(\nand_61.nand_4 )
  );
  nand2 \nand_61.nand2_5  (    .in_0(\nand_61.and_4 ),    .in_1(enable),    .out(\nand_61.out )
  );
  inverter \nand_62.inv_0  (    .in(\nand_62.nand_0 ),    .out(\nand_62.and_0 )
  );
  inverter \nand_62.inv_1  (    .in(\nand_62.nand_1 ),    .out(\nand_62.and_1 )
  );
  inverter \nand_62.inv_2  (    .in(\nand_62.nand_2 ),    .out(\nand_62.and_2 )
  );
  inverter \nand_62.inv_3  (    .in(\nand_62.nand_3 ),    .out(\nand_62.and_3 )
  );
  inverter \nand_62.inv_4  (    .in(\nand_62.nand_4 ),    .out(\nand_62.and_4 )
  );
  nand2 \nand_62.nand2_0  (    .in_0(\in_b<0> ),    .in_1(\in<1> ),    .out(\nand_62.nand_0 )
  );
  nand2 \nand_62.nand2_1  (    .in_0(\nand_62.and_0 ),    .in_1(\in<2> ),    .out(\nand_62.nand_1 )
  );
  nand2 \nand_62.nand2_2  (    .in_0(\nand_62.and_1 ),    .in_1(\in<3> ),    .out(\nand_62.nand_2 )
  );
  nand2 \nand_62.nand2_3  (    .in_0(\nand_62.and_2 ),    .in_1(\in<4> ),    .out(\nand_62.nand_3 )
  );
  nand2 \nand_62.nand2_4  (    .in_0(\nand_62.and_3 ),    .in_1(\in<5> ),    .out(\nand_62.nand_4 )
  );
  nand2 \nand_62.nand2_5  (    .in_0(\nand_62.and_4 ),    .in_1(enable),    .out(\nand_62.out )
  );
  inverter \nand_63.inv_0  (    .in(\nand_63.nand_0 ),    .out(\nand_63.and_0 )
  );
  inverter \nand_63.inv_1  (    .in(\nand_63.nand_1 ),    .out(\nand_63.and_1 )
  );
  inverter \nand_63.inv_2  (    .in(\nand_63.nand_2 ),    .out(\nand_63.and_2 )
  );
  inverter \nand_63.inv_3  (    .in(\nand_63.nand_3 ),    .out(\nand_63.and_3 )
  );
  inverter \nand_63.inv_4  (    .in(\nand_63.nand_4 ),    .out(\nand_63.and_4 )
  );
  nand2 \nand_63.nand2_0  (    .in_0(\in<0> ),    .in_1(\in<1> ),    .out(\nand_63.nand_0 )
  );
  nand2 \nand_63.nand2_1  (    .in_0(\nand_63.and_0 ),    .in_1(\in<2> ),    .out(\nand_63.nand_1 )
  );
  nand2 \nand_63.nand2_2  (    .in_0(\nand_63.and_1 ),    .in_1(\in<3> ),    .out(\nand_63.nand_2 )
  );
  nand2 \nand_63.nand2_3  (    .in_0(\nand_63.and_2 ),    .in_1(\in<4> ),    .out(\nand_63.nand_3 )
  );
  nand2 \nand_63.nand2_4  (    .in_0(\nand_63.and_3 ),    .in_1(\in<5> ),    .out(\nand_63.nand_4 )
  );
  nand2 \nand_63.nand2_5  (    .in_0(\nand_63.and_4 ),    .in_1(enable),    .out(\nand_63.out )
  );
  inverter \nand_7.inv_0  (    .in(\nand_7.nand_0 ),    .out(\nand_7.and_0 )
  );
  inverter \nand_7.inv_1  (    .in(\nand_7.nand_1 ),    .out(\nand_7.and_1 )
  );
  inverter \nand_7.inv_2  (    .in(\nand_7.nand_2 ),    .out(\nand_7.and_2 )
  );
  inverter \nand_7.inv_3  (    .in(\nand_7.nand_3 ),    .out(\nand_7.and_3 )
  );
  inverter \nand_7.inv_4  (    .in(\nand_7.nand_4 ),    .out(\nand_7.and_4 )
  );
  nand2 \nand_7.nand2_0  (    .in_0(\in<0> ),    .in_1(\in<1> ),    .out(\nand_7.nand_0 )
  );
  nand2 \nand_7.nand2_1  (    .in_0(\nand_7.and_0 ),    .in_1(\in<2> ),    .out(\nand_7.nand_1 )
  );
  nand2 \nand_7.nand2_2  (    .in_0(\nand_7.and_1 ),    .in_1(\in_b<3> ),    .out(\nand_7.nand_2 )
  );
  nand2 \nand_7.nand2_3  (    .in_0(\nand_7.and_2 ),    .in_1(\in_b<4> ),    .out(\nand_7.nand_3 )
  );
  nand2 \nand_7.nand2_4  (    .in_0(\nand_7.and_3 ),    .in_1(\in_b<5> ),    .out(\nand_7.nand_4 )
  );
  nand2 \nand_7.nand2_5  (    .in_0(\nand_7.and_4 ),    .in_1(enable),    .out(\nand_7.out )
  );
  inverter \nand_8.inv_0  (    .in(\nand_8.nand_0 ),    .out(\nand_8.and_0 )
  );
  inverter \nand_8.inv_1  (    .in(\nand_8.nand_1 ),    .out(\nand_8.and_1 )
  );
  inverter \nand_8.inv_2  (    .in(\nand_8.nand_2 ),    .out(\nand_8.and_2 )
  );
  inverter \nand_8.inv_3  (    .in(\nand_8.nand_3 ),    .out(\nand_8.and_3 )
  );
  inverter \nand_8.inv_4  (    .in(\nand_8.nand_4 ),    .out(\nand_8.and_4 )
  );
  nand2 \nand_8.nand2_0  (    .in_0(\in_b<0> ),    .in_1(\in_b<1> ),    .out(\nand_8.nand_0 )
  );
  nand2 \nand_8.nand2_1  (    .in_0(\nand_8.and_0 ),    .in_1(\in_b<2> ),    .out(\nand_8.nand_1 )
  );
  nand2 \nand_8.nand2_2  (    .in_0(\nand_8.and_1 ),    .in_1(\in<3> ),    .out(\nand_8.nand_2 )
  );
  nand2 \nand_8.nand2_3  (    .in_0(\nand_8.and_2 ),    .in_1(\in_b<4> ),    .out(\nand_8.nand_3 )
  );
  nand2 \nand_8.nand2_4  (    .in_0(\nand_8.and_3 ),    .in_1(\in_b<5> ),    .out(\nand_8.nand_4 )
  );
  nand2 \nand_8.nand2_5  (    .in_0(\nand_8.and_4 ),    .in_1(enable),    .out(\nand_8.out )
  );
  inverter \nand_9.inv_0  (    .in(\nand_9.nand_0 ),    .out(\nand_9.and_0 )
  );
  inverter \nand_9.inv_1  (    .in(\nand_9.nand_1 ),    .out(\nand_9.and_1 )
  );
  inverter \nand_9.inv_2  (    .in(\nand_9.nand_2 ),    .out(\nand_9.and_2 )
  );
  inverter \nand_9.inv_3  (    .in(\nand_9.nand_3 ),    .out(\nand_9.and_3 )
  );
  inverter \nand_9.inv_4  (    .in(\nand_9.nand_4 ),    .out(\nand_9.and_4 )
  );
  nand2 \nand_9.nand2_0  (    .in_0(\in<0> ),    .in_1(\in_b<1> ),    .out(\nand_9.nand_0 )
  );
  nand2 \nand_9.nand2_1  (    .in_0(\nand_9.and_0 ),    .in_1(\in_b<2> ),    .out(\nand_9.nand_1 )
  );
  nand2 \nand_9.nand2_2  (    .in_0(\nand_9.and_1 ),    .in_1(\in<3> ),    .out(\nand_9.nand_2 )
  );
  nand2 \nand_9.nand2_3  (    .in_0(\nand_9.and_2 ),    .in_1(\in_b<4> ),    .out(\nand_9.nand_3 )
  );
  nand2 \nand_9.nand2_4  (    .in_0(\nand_9.and_3 ),    .in_1(\in_b<5> ),    .out(\nand_9.nand_4 )
  );
  nand2 \nand_9.nand2_5  (    .in_0(\nand_9.and_4 ),    .in_1(enable),    .out(\nand_9.out )
  );
  assign \out_b<59>  = \nand_59.out ;
  assign \out_b<58>  = \nand_58.out ;
  assign \out_b<57>  = \nand_57.out ;
  assign \out_b<56>  = \nand_56.out ;
  assign \out_b<55>  = \nand_55.out ;
  assign \out_b<54>  = \nand_54.out ;
  assign \out_b<53>  = \nand_53.out ;
  assign \out_b<52>  = \nand_52.out ;
  assign \out_b<51>  = \nand_51.out ;
  assign \out_b<50>  = \nand_50.out ;
  assign \out_b<49>  = \nand_49.out ;
  assign \out_b<48>  = \nand_48.out ;
  assign \out_b<47>  = \nand_47.out ;
  assign \out_b<46>  = \nand_46.out ;
  assign \out_b<45>  = \nand_45.out ;
  assign \out_b<44>  = \nand_44.out ;
  assign \out_b<43>  = \nand_43.out ;
  assign \out_b<42>  = \nand_42.out ;
  assign \out_b<41>  = \nand_41.out ;
  assign \out_b<40>  = \nand_40.out ;
  assign \out_b<39>  = \nand_39.out ;
  assign \out_b<38>  = \nand_38.out ;
  assign \out_b<37>  = \nand_37.out ;
  assign \out_b<36>  = \nand_36.out ;
  assign \out_b<35>  = \nand_35.out ;
  assign \out_b<34>  = \nand_34.out ;
  assign \out_b<33>  = \nand_33.out ;
  assign \out_b<32>  = \nand_32.out ;
  assign \out_b<31>  = \nand_31.out ;
  assign \out_b<30>  = \nand_30.out ;
  assign \out_b<29>  = \nand_29.out ;
  assign \out_b<28>  = \nand_28.out ;
  assign \out_b<27>  = \nand_27.out ;
  assign \out_b<26>  = \nand_26.out ;
  assign \out_b<25>  = \nand_25.out ;
  assign \out_b<24>  = \nand_24.out ;
  assign \out_b<23>  = \nand_23.out ;
  assign \out_b<22>  = \nand_22.out ;
  assign \out_b<21>  = \nand_21.out ;
  assign \out_b<20>  = \nand_20.out ;
  assign \out_b<19>  = \nand_19.out ;
  assign \out_b<18>  = \nand_18.out ;
  assign \out_b<17>  = \nand_17.out ;
  assign \out_b<16>  = \nand_16.out ;
  assign \out_b<15>  = \nand_15.out ;
  assign \out_b<14>  = \nand_14.out ;
  assign \out_b<13>  = \nand_13.out ;
  assign \out_b<12>  = \nand_12.out ;
  assign \out_b<11>  = \nand_11.out ;
  assign \out_b<10>  = \nand_10.out ;
  assign \out_b<9>  = \nand_9.out ;
  assign \out_b<8>  = \nand_8.out ;
  assign \out_b<7>  = \nand_7.out ;
  assign \out_b<6>  = \nand_6.out ;
  assign \out_b<5>  = \nand_5.out ;
  assign \out_b<4>  = \nand_4.out ;
  assign \out_b<3>  = \nand_3.out ;
  assign \out_b<2>  = \nand_2.out ;
  assign \out_b<1>  = \nand_1.out ;
  assign \out_b<0>  = \nand_0.out ;
  assign \nand_63.in_0  = \in<0> ;
  assign \nand_63.in_1  = \in<1> ;
  assign \nand_63.in_2  = \in<2> ;
  assign \nand_63.in_3  = \in<3> ;
  assign \nand_63.in_4  = \in<4> ;
  assign \nand_63.in_5  = \in<5> ;
  assign \nand_63.in_6  = enable;
  assign \nand_62.in_0  = \in_b<0> ;
  assign \nand_62.in_1  = \in<1> ;
  assign \nand_62.in_2  = \in<2> ;
  assign \nand_62.in_3  = \in<3> ;
  assign \nand_62.in_4  = \in<4> ;
  assign \nand_62.in_5  = \in<5> ;
  assign \nand_62.in_6  = enable;
  assign \nand_61.in_0  = \in<0> ;
  assign \nand_61.in_1  = \in_b<1> ;
  assign \nand_61.in_2  = \in<2> ;
  assign \nand_61.in_3  = \in<3> ;
  assign \nand_61.in_4  = \in<4> ;
  assign \nand_61.in_5  = \in<5> ;
  assign \nand_61.in_6  = enable;
  assign \nand_60.in_0  = \in_b<0> ;
  assign \nand_60.in_1  = \in_b<1> ;
  assign \nand_60.in_2  = \in<2> ;
  assign \nand_60.in_3  = \in<3> ;
  assign \nand_60.in_4  = \in<4> ;
  assign \nand_60.in_5  = \in<5> ;
  assign \nand_60.in_6  = enable;
  assign \nand_59.in_0  = \in<0> ;
  assign \nand_59.in_1  = \in<1> ;
  assign \nand_59.in_2  = \in_b<2> ;
  assign \nand_59.in_3  = \in<3> ;
  assign \nand_59.in_4  = \in<4> ;
  assign \nand_59.in_5  = \in<5> ;
  assign \nand_59.in_6  = enable;
  assign \nand_58.in_0  = \in_b<0> ;
  assign \nand_58.in_1  = \in<1> ;
  assign \nand_58.in_2  = \in_b<2> ;
  assign \nand_58.in_3  = \in<3> ;
  assign \nand_58.in_4  = \in<4> ;
  assign \nand_58.in_5  = \in<5> ;
  assign \nand_58.in_6  = enable;
  assign \nand_57.in_0  = \in<0> ;
  assign \nand_57.in_1  = \in_b<1> ;
  assign \nand_57.in_2  = \in_b<2> ;
  assign \nand_57.in_3  = \in<3> ;
  assign \nand_57.in_4  = \in<4> ;
  assign \nand_57.in_5  = \in<5> ;
  assign \nand_57.in_6  = enable;
  assign \nand_56.in_0  = \in_b<0> ;
  assign \nand_56.in_1  = \in_b<1> ;
  assign \nand_56.in_2  = \in_b<2> ;
  assign \nand_56.in_3  = \in<3> ;
  assign \nand_56.in_4  = \in<4> ;
  assign \nand_56.in_5  = \in<5> ;
  assign \nand_56.in_6  = enable;
  assign \nand_55.in_0  = \in<0> ;
  assign \nand_55.in_1  = \in<1> ;
  assign \nand_55.in_2  = \in<2> ;
  assign \nand_55.in_3  = \in_b<3> ;
  assign \nand_55.in_4  = \in<4> ;
  assign \nand_55.in_5  = \in<5> ;
  assign \nand_55.in_6  = enable;
  assign \nand_54.in_0  = \in_b<0> ;
  assign \nand_54.in_1  = \in<1> ;
  assign \nand_54.in_2  = \in<2> ;
  assign \nand_54.in_3  = \in_b<3> ;
  assign \nand_54.in_4  = \in<4> ;
  assign \nand_54.in_5  = \in<5> ;
  assign \nand_54.in_6  = enable;
  assign \nand_53.in_0  = \in<0> ;
  assign \nand_53.in_1  = \in_b<1> ;
  assign \nand_53.in_2  = \in<2> ;
  assign \nand_53.in_3  = \in_b<3> ;
  assign \nand_53.in_4  = \in<4> ;
  assign \nand_53.in_5  = \in<5> ;
  assign \nand_53.in_6  = enable;
  assign \nand_52.in_0  = \in_b<0> ;
  assign \nand_52.in_1  = \in_b<1> ;
  assign \nand_52.in_2  = \in<2> ;
  assign \nand_52.in_3  = \in_b<3> ;
  assign \nand_52.in_4  = \in<4> ;
  assign \nand_52.in_5  = \in<5> ;
  assign \nand_52.in_6  = enable;
  assign \nand_51.in_0  = \in<0> ;
  assign \nand_51.in_1  = \in<1> ;
  assign \nand_51.in_2  = \in_b<2> ;
  assign \nand_51.in_3  = \in_b<3> ;
  assign \nand_51.in_4  = \in<4> ;
  assign \nand_51.in_5  = \in<5> ;
  assign \nand_51.in_6  = enable;
  assign \nand_50.in_0  = \in_b<0> ;
  assign \nand_50.in_1  = \in<1> ;
  assign \nand_50.in_2  = \in_b<2> ;
  assign \nand_50.in_3  = \in_b<3> ;
  assign \nand_50.in_4  = \in<4> ;
  assign \nand_50.in_5  = \in<5> ;
  assign \nand_50.in_6  = enable;
  assign \nand_49.in_0  = \in<0> ;
  assign \nand_49.in_1  = \in_b<1> ;
  assign \nand_49.in_2  = \in_b<2> ;
  assign \nand_49.in_3  = \in_b<3> ;
  assign \nand_49.in_4  = \in<4> ;
  assign \nand_49.in_5  = \in<5> ;
  assign \nand_49.in_6  = enable;
  assign \nand_48.in_0  = \in_b<0> ;
  assign \nand_48.in_1  = \in_b<1> ;
  assign \nand_48.in_2  = \in_b<2> ;
  assign \nand_48.in_3  = \in_b<3> ;
  assign \nand_48.in_4  = \in<4> ;
  assign \nand_48.in_5  = \in<5> ;
  assign \nand_48.in_6  = enable;
  assign \nand_47.in_0  = \in<0> ;
  assign \nand_47.in_1  = \in<1> ;
  assign \nand_47.in_2  = \in<2> ;
  assign \nand_47.in_3  = \in<3> ;
  assign \nand_47.in_4  = \in_b<4> ;
  assign \nand_47.in_5  = \in<5> ;
  assign \nand_47.in_6  = enable;
  assign \nand_46.in_0  = \in_b<0> ;
  assign \nand_46.in_1  = \in<1> ;
  assign \nand_46.in_2  = \in<2> ;
  assign \nand_46.in_3  = \in<3> ;
  assign \nand_46.in_4  = \in_b<4> ;
  assign \nand_46.in_5  = \in<5> ;
  assign \nand_46.in_6  = enable;
  assign \nand_45.in_0  = \in<0> ;
  assign \nand_45.in_1  = \in_b<1> ;
  assign \nand_45.in_2  = \in<2> ;
  assign \nand_45.in_3  = \in<3> ;
  assign \nand_45.in_4  = \in_b<4> ;
  assign \nand_45.in_5  = \in<5> ;
  assign \nand_45.in_6  = enable;
  assign \nand_44.in_0  = \in_b<0> ;
  assign \nand_44.in_1  = \in_b<1> ;
  assign \nand_44.in_2  = \in<2> ;
  assign \nand_44.in_3  = \in<3> ;
  assign \nand_44.in_4  = \in_b<4> ;
  assign \nand_44.in_5  = \in<5> ;
  assign \nand_44.in_6  = enable;
  assign \nand_43.in_0  = \in<0> ;
  assign \nand_43.in_1  = \in<1> ;
  assign \nand_43.in_2  = \in_b<2> ;
  assign \nand_43.in_3  = \in<3> ;
  assign \nand_43.in_4  = \in_b<4> ;
  assign \nand_43.in_5  = \in<5> ;
  assign \nand_43.in_6  = enable;
  assign \nand_42.in_0  = \in_b<0> ;
  assign \nand_42.in_1  = \in<1> ;
  assign \nand_42.in_2  = \in_b<2> ;
  assign \nand_42.in_3  = \in<3> ;
  assign \nand_42.in_4  = \in_b<4> ;
  assign \nand_42.in_5  = \in<5> ;
  assign \nand_42.in_6  = enable;
  assign \nand_41.in_0  = \in<0> ;
  assign \nand_41.in_1  = \in_b<1> ;
  assign \nand_41.in_2  = \in_b<2> ;
  assign \nand_41.in_3  = \in<3> ;
  assign \nand_41.in_4  = \in_b<4> ;
  assign \nand_41.in_5  = \in<5> ;
  assign \nand_41.in_6  = enable;
  assign \nand_40.in_0  = \in_b<0> ;
  assign \nand_40.in_1  = \in_b<1> ;
  assign \nand_40.in_2  = \in_b<2> ;
  assign \nand_40.in_3  = \in<3> ;
  assign \nand_40.in_4  = \in_b<4> ;
  assign \nand_40.in_5  = \in<5> ;
  assign \nand_40.in_6  = enable;
  assign \nand_39.in_0  = \in<0> ;
  assign \nand_39.in_1  = \in<1> ;
  assign \nand_39.in_2  = \in<2> ;
  assign \nand_39.in_3  = \in_b<3> ;
  assign \nand_39.in_4  = \in_b<4> ;
  assign \nand_39.in_5  = \in<5> ;
  assign \nand_39.in_6  = enable;
  assign \nand_38.in_0  = \in_b<0> ;
  assign \nand_38.in_1  = \in<1> ;
  assign \nand_38.in_2  = \in<2> ;
  assign \nand_38.in_3  = \in_b<3> ;
  assign \nand_38.in_4  = \in_b<4> ;
  assign \nand_38.in_5  = \in<5> ;
  assign \nand_38.in_6  = enable;
  assign \nand_37.in_0  = \in<0> ;
  assign \nand_37.in_1  = \in_b<1> ;
  assign \nand_37.in_2  = \in<2> ;
  assign \nand_37.in_3  = \in_b<3> ;
  assign \nand_37.in_4  = \in_b<4> ;
  assign \nand_37.in_5  = \in<5> ;
  assign \nand_37.in_6  = enable;
  assign \nand_36.in_0  = \in_b<0> ;
  assign \nand_36.in_1  = \in_b<1> ;
  assign \nand_36.in_2  = \in<2> ;
  assign \nand_36.in_3  = \in_b<3> ;
  assign \nand_36.in_4  = \in_b<4> ;
  assign \nand_36.in_5  = \in<5> ;
  assign \nand_36.in_6  = enable;
  assign \nand_35.in_0  = \in<0> ;
  assign \nand_35.in_1  = \in<1> ;
  assign \nand_35.in_2  = \in_b<2> ;
  assign \nand_35.in_3  = \in_b<3> ;
  assign \nand_35.in_4  = \in_b<4> ;
  assign \nand_35.in_5  = \in<5> ;
  assign \nand_35.in_6  = enable;
  assign \nand_34.in_0  = \in_b<0> ;
  assign \nand_34.in_1  = \in<1> ;
  assign \nand_34.in_2  = \in_b<2> ;
  assign \nand_34.in_3  = \in_b<3> ;
  assign \nand_34.in_4  = \in_b<4> ;
  assign \nand_34.in_5  = \in<5> ;
  assign \nand_34.in_6  = enable;
  assign \nand_33.in_0  = \in<0> ;
  assign \nand_33.in_1  = \in_b<1> ;
  assign \nand_33.in_2  = \in_b<2> ;
  assign \nand_33.in_3  = \in_b<3> ;
  assign \nand_33.in_4  = \in_b<4> ;
  assign \nand_33.in_5  = \in<5> ;
  assign \nand_33.in_6  = enable;
  assign \nand_32.in_0  = \in_b<0> ;
  assign \nand_32.in_1  = \in_b<1> ;
  assign \nand_32.in_2  = \in_b<2> ;
  assign \nand_32.in_3  = \in_b<3> ;
  assign \nand_32.in_4  = \in_b<4> ;
  assign \nand_32.in_5  = \in<5> ;
  assign \nand_32.in_6  = enable;
  assign \nand_31.in_0  = \in<0> ;
  assign \nand_31.in_1  = \in<1> ;
  assign \nand_31.in_2  = \in<2> ;
  assign \nand_31.in_3  = \in<3> ;
  assign \nand_31.in_4  = \in<4> ;
  assign \nand_31.in_5  = \in_b<5> ;
  assign \nand_31.in_6  = enable;
  assign \nand_30.in_0  = \in_b<0> ;
  assign \nand_30.in_1  = \in<1> ;
  assign \nand_30.in_2  = \in<2> ;
  assign \nand_30.in_3  = \in<3> ;
  assign \nand_30.in_4  = \in<4> ;
  assign \nand_30.in_5  = \in_b<5> ;
  assign \nand_30.in_6  = enable;
  assign \nand_29.in_0  = \in<0> ;
  assign \nand_29.in_1  = \in_b<1> ;
  assign \nand_29.in_2  = \in<2> ;
  assign \nand_29.in_3  = \in<3> ;
  assign \nand_29.in_4  = \in<4> ;
  assign \nand_29.in_5  = \in_b<5> ;
  assign \nand_29.in_6  = enable;
  assign \nand_28.in_0  = \in_b<0> ;
  assign \nand_28.in_1  = \in_b<1> ;
  assign \nand_28.in_2  = \in<2> ;
  assign \nand_28.in_3  = \in<3> ;
  assign \nand_28.in_4  = \in<4> ;
  assign \nand_28.in_5  = \in_b<5> ;
  assign \nand_28.in_6  = enable;
  assign \nand_27.in_0  = \in<0> ;
  assign \nand_27.in_1  = \in<1> ;
  assign \nand_27.in_2  = \in_b<2> ;
  assign \nand_27.in_3  = \in<3> ;
  assign \nand_27.in_4  = \in<4> ;
  assign \nand_27.in_5  = \in_b<5> ;
  assign \nand_27.in_6  = enable;
  assign \nand_26.in_0  = \in_b<0> ;
  assign \nand_26.in_1  = \in<1> ;
  assign \nand_26.in_2  = \in_b<2> ;
  assign \nand_26.in_3  = \in<3> ;
  assign \nand_26.in_4  = \in<4> ;
  assign \nand_26.in_5  = \in_b<5> ;
  assign \nand_26.in_6  = enable;
  assign \nand_25.in_0  = \in<0> ;
  assign \nand_25.in_1  = \in_b<1> ;
  assign \nand_25.in_2  = \in_b<2> ;
  assign \nand_25.in_3  = \in<3> ;
  assign \nand_25.in_4  = \in<4> ;
  assign \nand_25.in_5  = \in_b<5> ;
  assign \nand_25.in_6  = enable;
  assign \nand_24.in_0  = \in_b<0> ;
  assign \nand_24.in_1  = \in_b<1> ;
  assign \nand_24.in_2  = \in_b<2> ;
  assign \nand_24.in_3  = \in<3> ;
  assign \nand_24.in_4  = \in<4> ;
  assign \nand_24.in_5  = \in_b<5> ;
  assign \nand_24.in_6  = enable;
  assign \nand_23.in_0  = \in<0> ;
  assign \nand_23.in_1  = \in<1> ;
  assign \nand_23.in_2  = \in<2> ;
  assign \nand_23.in_3  = \in_b<3> ;
  assign \nand_23.in_4  = \in<4> ;
  assign \nand_23.in_5  = \in_b<5> ;
  assign \nand_23.in_6  = enable;
  assign \nand_22.in_0  = \in_b<0> ;
  assign \nand_22.in_1  = \in<1> ;
  assign \nand_22.in_2  = \in<2> ;
  assign \nand_22.in_3  = \in_b<3> ;
  assign \nand_22.in_4  = \in<4> ;
  assign \nand_22.in_5  = \in_b<5> ;
  assign \nand_22.in_6  = enable;
  assign \nand_21.in_0  = \in<0> ;
  assign \nand_21.in_1  = \in_b<1> ;
  assign \nand_21.in_2  = \in<2> ;
  assign \nand_21.in_3  = \in_b<3> ;
  assign \nand_21.in_4  = \in<4> ;
  assign \nand_21.in_5  = \in_b<5> ;
  assign \nand_21.in_6  = enable;
  assign \nand_20.in_0  = \in_b<0> ;
  assign \nand_20.in_1  = \in_b<1> ;
  assign \nand_20.in_2  = \in<2> ;
  assign \nand_20.in_3  = \in_b<3> ;
  assign \nand_20.in_4  = \in<4> ;
  assign \nand_20.in_5  = \in_b<5> ;
  assign \nand_20.in_6  = enable;
  assign \nand_19.in_0  = \in<0> ;
  assign \nand_19.in_1  = \in<1> ;
  assign \nand_19.in_2  = \in_b<2> ;
  assign \nand_19.in_3  = \in_b<3> ;
  assign \nand_19.in_4  = \in<4> ;
  assign \nand_19.in_5  = \in_b<5> ;
  assign \nand_19.in_6  = enable;
  assign \nand_18.in_0  = \in_b<0> ;
  assign \nand_18.in_1  = \in<1> ;
  assign \nand_18.in_2  = \in_b<2> ;
  assign \nand_18.in_3  = \in_b<3> ;
  assign \nand_18.in_4  = \in<4> ;
  assign \nand_18.in_5  = \in_b<5> ;
  assign \nand_18.in_6  = enable;
  assign \nand_17.in_0  = \in<0> ;
  assign \nand_17.in_1  = \in_b<1> ;
  assign \nand_17.in_2  = \in_b<2> ;
  assign \nand_17.in_3  = \in_b<3> ;
  assign \nand_17.in_4  = \in<4> ;
  assign \nand_17.in_5  = \in_b<5> ;
  assign \nand_17.in_6  = enable;
  assign \nand_16.in_0  = \in_b<0> ;
  assign \nand_16.in_1  = \in_b<1> ;
  assign \nand_16.in_2  = \in_b<2> ;
  assign \nand_16.in_3  = \in_b<3> ;
  assign \nand_16.in_4  = \in<4> ;
  assign \nand_16.in_5  = \in_b<5> ;
  assign \nand_16.in_6  = enable;
  assign \nand_15.in_0  = \in<0> ;
  assign \nand_15.in_1  = \in<1> ;
  assign \nand_15.in_2  = \in<2> ;
  assign \nand_15.in_3  = \in<3> ;
  assign \nand_15.in_4  = \in_b<4> ;
  assign \nand_15.in_5  = \in_b<5> ;
  assign \nand_15.in_6  = enable;
  assign \nand_14.in_0  = \in_b<0> ;
  assign \nand_14.in_1  = \in<1> ;
  assign \nand_14.in_2  = \in<2> ;
  assign \nand_14.in_3  = \in<3> ;
  assign \nand_14.in_4  = \in_b<4> ;
  assign \nand_14.in_5  = \in_b<5> ;
  assign \nand_14.in_6  = enable;
  assign \nand_13.in_0  = \in<0> ;
  assign \nand_13.in_1  = \in_b<1> ;
  assign \nand_13.in_2  = \in<2> ;
  assign \nand_13.in_3  = \in<3> ;
  assign \nand_13.in_4  = \in_b<4> ;
  assign \nand_13.in_5  = \in_b<5> ;
  assign \nand_13.in_6  = enable;
  assign \nand_12.in_0  = \in_b<0> ;
  assign \nand_12.in_1  = \in_b<1> ;
  assign \nand_12.in_2  = \in<2> ;
  assign \nand_12.in_3  = \in<3> ;
  assign \nand_12.in_4  = \in_b<4> ;
  assign \nand_12.in_5  = \in_b<5> ;
  assign \nand_12.in_6  = enable;
  assign \nand_11.in_0  = \in<0> ;
  assign \nand_11.in_1  = \in<1> ;
  assign \nand_11.in_2  = \in_b<2> ;
  assign \nand_11.in_3  = \in<3> ;
  assign \nand_11.in_4  = \in_b<4> ;
  assign \nand_11.in_5  = \in_b<5> ;
  assign \nand_11.in_6  = enable;
  assign \nand_10.in_0  = \in_b<0> ;
  assign \nand_10.in_1  = \in<1> ;
  assign \nand_10.in_2  = \in_b<2> ;
  assign \nand_10.in_3  = \in<3> ;
  assign \nand_10.in_4  = \in_b<4> ;
  assign \nand_10.in_5  = \in_b<5> ;
  assign \nand_10.in_6  = enable;
  assign \nand_9.in_0  = \in<0> ;
  assign \nand_9.in_1  = \in_b<1> ;
  assign \nand_9.in_2  = \in_b<2> ;
  assign \nand_9.in_3  = \in<3> ;
  assign \nand_9.in_4  = \in_b<4> ;
  assign \nand_9.in_5  = \in_b<5> ;
  assign \nand_9.in_6  = enable;
  assign \nand_8.in_0  = \in_b<0> ;
  assign \nand_8.in_1  = \in_b<1> ;
  assign \nand_8.in_2  = \in_b<2> ;
  assign \nand_8.in_3  = \in<3> ;
  assign \nand_8.in_4  = \in_b<4> ;
  assign \nand_8.in_5  = \in_b<5> ;
  assign \nand_8.in_6  = enable;
  assign \nand_7.in_0  = \in<0> ;
  assign \nand_7.in_1  = \in<1> ;
  assign \nand_7.in_2  = \in<2> ;
  assign \nand_7.in_3  = \in_b<3> ;
  assign \nand_7.in_4  = \in_b<4> ;
  assign \nand_7.in_5  = \in_b<5> ;
  assign \nand_7.in_6  = enable;
  assign \nand_6.in_0  = \in_b<0> ;
  assign \nand_6.in_1  = \in<1> ;
  assign \nand_6.in_2  = \in<2> ;
  assign \nand_6.in_3  = \in_b<3> ;
  assign \nand_6.in_4  = \in_b<4> ;
  assign \nand_6.in_5  = \in_b<5> ;
  assign \nand_6.in_6  = enable;
  assign \nand_5.in_0  = \in<0> ;
  assign \nand_5.in_1  = \in_b<1> ;
  assign \nand_5.in_2  = \in<2> ;
  assign \nand_5.in_3  = \in_b<3> ;
  assign \nand_5.in_4  = \in_b<4> ;
  assign \nand_5.in_5  = \in_b<5> ;
  assign \nand_5.in_6  = enable;
  assign \nand_4.in_0  = \in_b<0> ;
  assign \nand_4.in_1  = \in_b<1> ;
  assign \nand_4.in_2  = \in<2> ;
  assign \nand_4.in_3  = \in_b<3> ;
  assign \nand_4.in_4  = \in_b<4> ;
  assign \nand_4.in_5  = \in_b<5> ;
  assign \nand_4.in_6  = enable;
  assign \nand_3.in_0  = \in<0> ;
  assign \nand_3.in_1  = \in<1> ;
  assign \nand_3.in_2  = \in_b<2> ;
  assign \nand_3.in_3  = \in_b<3> ;
  assign \nand_3.in_4  = \in_b<4> ;
  assign \nand_3.in_5  = \in_b<5> ;
  assign \nand_3.in_6  = enable;
  assign \nand_2.in_0  = \in_b<0> ;
  assign \nand_2.in_1  = \in<1> ;
  assign \nand_2.in_2  = \in_b<2> ;
  assign \nand_2.in_3  = \in_b<3> ;
  assign \nand_2.in_4  = \in_b<4> ;
  assign \nand_2.in_5  = \in_b<5> ;
  assign \nand_2.in_6  = enable;
  assign \nand_1.in_0  = \in<0> ;
  assign \nand_1.in_1  = \in_b<1> ;
  assign \nand_1.in_2  = \in_b<2> ;
  assign \nand_1.in_3  = \in_b<3> ;
  assign \nand_1.in_4  = \in_b<4> ;
  assign \nand_1.in_5  = \in_b<5> ;
  assign \nand_1.in_6  = enable;
  assign \nand_0.in_0  = \in_b<0> ;
  assign \nand_0.in_1  = \in_b<1> ;
  assign \nand_0.in_2  = \in_b<2> ;
  assign \nand_0.in_3  = \in_b<3> ;
  assign \nand_0.in_4  = \in_b<4> ;
  assign \nand_0.in_5  = \in_b<5> ;
  assign \nand_0.in_6  = enable;
  assign \out_b<63>  = \nand_63.out ;
  assign \out_b<62>  = \nand_62.out ;
  assign \out_b<61>  = \nand_61.out ;
  assign \out_b<60>  = \nand_60.out ;
endmodule
